--
-- Simplistic 4096x16 rom module
--
-- This source code is public domain
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
port (
   CLK  : in  std_logic;
   nCS  : in  std_logic;
   ADDR : in  std_logic_vector (11 downto 0);    -- note: word adress!
   DO   : out std_logic_vector (15 downto 0)
   );
end rom;

--ROM content: Stuart's EVMBUG rom, first 8KB

architecture rom_arch of rom is

   constant size : integer := 4095;
	type mem_array is array(0 to size) of std_logic_vector(15 downto 0);
	constant rom : mem_array := (                                              -- byte addr:
		x"ec00", x"0226", x"f0d6", x"f0f6", x"f0ca", x"f0ea", x"f0be", x"f0de", -- address 0x0000
		x"f0b2", x"f0d2", x"0d0a", x"4d4f", x"4e3f", x"2000", x"2020", x"2020", -- address 0x0010
		x"2020", x"000d", x"0a42", x"5000", x"4944", x"543d", x"000d", x"0a52", -- address 0x0020
		x"4541", x"4459", x"2059", x"2f4e", x"2000", x"5700", x"5000", x"5300", -- address 0x0030
		x"f0ac", x"f0be", x"f09e", x"f0b0", x"f090", x"f0a2", x"f082", x"f094", -- address 0x0040
		x"f074", x"f086", x"f066", x"f078", x"f058", x"f06a", x"f04a", x"f05c", -- address 0x0050
		x"ec24", x"03f8", x"ec24", x"0396", x"ec24", x"0402", x"ec0a", x"0326", -- address 0x0060
		x"ec16", x"02ee", x"ec16", x"02e2", x"ec24", x"032c", x"ec00", x"0442", -- address 0x0070
		x"0460", x"0142", x"0009", x"0034", x"0012", x"0034", x"0023", x"0034", -- address 0x0080
		x"0046", x"0034", x"008d", x"0034", x"0119", x"0034", x"02a4", x"0034", -- address 0x0090
		x"7fff", x"0034", x"0d0a", x"4552", x"524f", x"5220", x"000d", x"0a45", -- address 0x00a0
		x"564d", x"4255", x"4720", x"2052", x"312e", x"3000", x"0d0a", x"5200", -- address 0x00b0
		x"0d0a", x"4831", x"2b48", x"323d", x"0020", x"4831", x"2d48", x"323d", -- address 0x00c0
		x"0020", x"4552", x"524f", x"5200", x"0d0a", x"434f", x"4d3f", x"2000", -- address 0x00d0
		x"3a0d", x"000d", x"0a54", x"4552", x"4d49", x"4e41", x"4c20", x"4d4f", -- address 0x00e0
		x"4445", x"0d0a", x"000d", x"0a43", x"4d44", x"2045", x"5252", x"000d", -- address 0x00f0
		x"0a50", x"4152", x"4d20", x"4552", x"5200", x"0d0a", x"434b", x"534d", -- address 0x0100
		x"2045", x"5252", x"000d", x"0a54", x"4147", x"2045", x"5252", x"0055", -- address 0x0110
		x"504c", x"4420", x"4552", x"5200", x"460d", x"000a", x"7f3a", x"0d0a", -- address 0x0120
		x"7f13", x"0d14", x"7f00", x"120a", x"7f00", x"6242", x"1100", x"0000", -- address 0x0130
		x"0400", x"02e0", x"ec00", x"04c1", x"0202", x"fffc", x"ccb1", x"0201", -- address 0x0140
		x"042e", x"cc81", x"0209", x"0142", x"04c1", x"0641", x"16fe", x"c320", -- address 0x0150
		x"013e", x"c80c", x"ec2e", x"1f15", x"1601", x"2f45", x"2fa0", x"0014", -- address 0x0160
		x"04c0", x"0202", x"0a05", x"0203", x"0004", x"04c4", x"0208", x"0001", -- address 0x0170
		x"2ec5", x"0285", x"0d00", x"1604", x"0205", x"0a00", x"2f05", x"1019", -- address 0x0180
		x"0285", x"2000", x"1316", x"0285", x"2c00", x"1313", x"0285", x"4100", -- address 0x0190
		x"113c", x"0285", x"5a00", x"1539", x"0603", x"1337", x"06c5", x"0245", -- address 0x01a0
		x"001f", x"0283", x"0003", x"1301", x"0482", x"a105", x"0222", x"0050", -- address 0x01b0
		x"10df", x"020b", x"027a", x"1002", x"022b", x"0004", x"c2bb", x"1325", -- address 0x01c0
		x"810a", x"16fa", x"c1bb", x"c2db", x"0207", x"ec00", x"0285", x"0a00", -- address 0x01d0
		x"130f", x"0916", x"170e", x"2e44", x"01f8", x"020e", x"cdc4", x"0583", -- address 0x01e0
		x"0285", x"0d00", x"1306", x"10f5", x"05c7", x"0285", x"0d00", x"16f7", -- address 0x01f0
		x"04c3", x"045b", x"04c0", x"100b", x"0200", x"0001", x"1008", x"0200", -- address 0x0200
		x"0002", x"1005", x"0200", x"0003", x"1002", x"0200", x"0004", x"2fa0", -- address 0x0210
		x"00a4", x"2e00", x"108e", x"020c", x"ec44", x"04fc", x"073c", x"04fc", -- address 0x0220
		x"04dc", x"c320", x"013e", x"c80c", x"ec2e", x"1d1f", x"04c3", x"3220", -- address 0x0230
		x"013a", x"1e0d", x"1f0f", x"13fe", x"0583", x"1f0f", x"16fd", x"0207", -- address 0x0240
		x"0084", x"8dc3", x"1102", x"05c7", x"10fc", x"3317", x"c1d7", x"0287", -- address 0x0250
		x"01a1", x"1108", x"1602", x"0720", x"ec44", x"2f45", x"2fa0", x"00ad", -- address 0x0260
		x"0460", x"0142", x"05a0", x"ec44", x"10f8", x"01a9", x"0001", x"036c", -- address 0x0270
		x"01a4", x"0003", x"0334", x"4ae9", x"0001", x"04ac", x"0305", x"0000", -- address 0x0280
		x"042c", x"0b05", x"0001", x"0436", x"0273", x"0000", x"0426", x"0dac", -- address 0x0290
		x"0001", x"064a", x"0da4", x"0007", x"0552", x"0069", x"0003", x"0460", -- address 0x02a0
		x"0249", x"0000", x"051a", x"0086", x"0007", x"0770", x"60a8", x"0003", -- address 0x02b0
		x"07a0", x"19d4", x"0000", x"07b4", x"1438", x"0001", x"07c2", x"0038", -- address 0x02c0
		x"0001", x"07ba", x"3078", x"0000", x"0e1a", x"0658", x"0003", x"1166", -- address 0x02d0
		x"0000", x"1f15", x"16fe", x"04db", x"361b", x"1e12", x"0380", x"020a", -- address 0x02e0
		x"186a", x"1d10", x"1f16", x"16fe", x"321b", x"d2db", x"980b", x"00f2", -- address 0x02f0
		x"160b", x"c2e0", x"ec44", x"150e", x"0a3a", x"1f16", x"16fe", x"1f17", -- address 0x0300
		x"16fc", x"060a", x"16fe", x"0380", x"c2e0", x"ec46", x"1303", x"c2e0", -- address 0x0310
		x"ec44", x"11f3", x"0380", x"2f5b", x"2f1b", x"0380", x"d33b", x"13fd", -- address 0x0320
		x"2f0c", x"10fc", x"4008", x"4048", x"0203", x"0008", x"2fa0", x"00f2", -- address 0x0330
		x"2e80", x"2fa0", x"00cf", x"2e90", x"1f15", x"1602", x"2f40", x"0459", -- address 0x0340
		x"8040", x"13fd", x"05c0", x"0603", x"0283", x"0004", x"1602", x"2fa0", -- address 0x0350
		x"0020", x"c0c3", x"13e9", x"2fa0", x"0020", x"10ed", x"4008", x"1004", -- address 0x0360
		x"0640", x"0a25", x"16fb", x"8c30", x"2fa0", x"00f2", x"2e80", x"2fa0", -- address 0x0370
		x"00cf", x"2e90", x"2fa0", x"0020", x"2e44", x"0390", x"020e", x"c404", -- address 0x0380
		x"0a25", x"11ee", x"0459", x"04c9", x"04cc", x"2eca", x"028a", x"3000", -- address 0x0390
		x"1a11", x"028a", x"3900", x"1208", x"028a", x"4100", x"1a0b", x"028a", -- address 0x03a0
		x"4600", x"1b08", x"022a", x"0900", x"0a4a", x"09ca", x"0a4c", x"a30a", -- address 0x03b0
		x"0589", x"10eb", x"028a", x"2000", x"130b", x"028a", x"2d00", x"1308", -- address 0x03c0
		x"028a", x"0d00", x"1305", x"028a", x"2c00", x"160c", x"020a", x"2000", -- address 0x03d0
		x"c249", x"1304", x"cecc", x"c6ca", x"8fbe", x"0380", x"05cb", x"c6ca", -- address 0x03e0
		x"c39e", x"0380", x"05ce", x"10fc", x"c31b", x"0acc", x"0209", x"0001", -- address 0x03f0
		x"1003", x"c31b", x"0209", x"0004", x"c28c", x"09ca", x"0a8a", x"028a", -- address 0x0400
		x"0900", x"1202", x"022a", x"0700", x"022a", x"3000", x"2f0a", x"0bcc", -- address 0x0410
		x"0609", x"16f2", x"0380", x"0207", x"9900", x"03e0", x"0380", x"0287", -- address 0x0420
		x"9900", x"130b", x"1013", x"4008", x"c190", x"c420", x"0440", x"0380", -- address 0x0430
		x"2fc0", x"064e", x"c406", x"2fa0", x"0023", x"04c7", x"020a", x"fffa", -- address 0x0440
		x"2fa0", x"001e", x"2eaa", x"ec20", x"05ca", x"16fa", x"0460", x"0142", -- address 0x0450
		x"c300", x"04c7", x"0241", x"000f", x"1303", x"0281", x"0009", x"1a01", -- address 0x0460
		x"0587", x"0a61", x"0208", x"3406", x"e201", x"0488", x"2fa0", x"00f2", -- address 0x0470
		x"2e8c", x"2fa0", x"00cf", x"c1c7", x"1601", x"0986", x"2e86", x"2fa0", -- address 0x0480
		x"0020", x"2e44", x"04a6", x"020e", x"c184", x"c1c7", x"1601", x"0a86", -- address 0x0490
		x"0248", x"f3ff", x"0488", x"09c5", x"16e5", x"0459", x"c1cd", x"c0c3", -- address 0x04a0
		x"131f", x"0240", x"000f", x"c180", x"0a10", x"a1c0", x"2fa0", x"00bc", -- address 0x04b0
		x"2e06", x"2fa0", x"00cf", x"2e97", x"2fa0", x"0020", x"2e44", x"04d4", -- address 0x04c0
		x"020e", x"c5c4", x"0a25", x"153c", x"0a15", x"1304", x"0606", x"1138", -- address 0x04d0
		x"0647", x"10ec", x"0286", x"000f", x"1333", x"0586", x"05c7", x"10e6", -- address 0x04e0
		x"04c6", x"c1cd", x"2fa0", x"00bc", x"2e06", x"2fa0", x"00cf", x"2e97", -- address 0x04f0
		x"0586", x"05c7", x"0286", x"0008", x"13f5", x"0286", x"0010", x"1320", -- address 0x0500
		x"2fa0", x"0020", x"2fa0", x"00d6", x"10ef", x"0206", x"003a", x"0207", -- address 0x0510
		x"0003", x"0208", x"ec1a", x"2fa0", x"00f2", x"2f96", x"2fa0", x"00cf", -- address 0x0520
		x"c118", x"2e98", x"2fa0", x"0020", x"2e44", x"053e", x"020e", x"c604", -- address 0x0530
		x"0a25", x"1506", x"0a15", x"16ef", x"05c6", x"05c8", x"0607", x"16eb", -- address 0x0540
		x"0459", x"4008", x"4048", x"4088", x"8040", x"1202", x"0460", x"0214", -- address 0x0550
		x"04c4", x"04c3", x"2fa0", x"0028", x"2f44", x"0284", x"0d00", x"1603", -- address 0x0560
		x"0204", x"2000", x"1001", x"2f04", x"d8c4", x"ec0c", x"0583", x"0283", -- address 0x0570
		x"0008", x"1304", x"0284", x"2000", x"16ef", x"10f6", x"2fa0", x"002d", -- address 0x0580
		x"2f44", x"0284", x"5900", x"1641", x"04e0", x"ec46", x"2fa0", x"0136", -- address 0x0590
		x"04ca", x"04c5", x"06a0", x"061c", x"3000", x"2fa0", x"ec0c", x"0203", -- address 0x05a0
		x"0008", x"d123", x"ec0b", x"0984", x"a144", x"0603", x"16fa", x"c282", -- address 0x05b0
		x"06a0", x"061c", x"3100", x"c280", x"06a0", x"061c", x"3900", x"c290", -- address 0x05c0
		x"06a0", x"061c", x"4200", x"8040", x"1304", x"05c0", x"0283", x"003c", -- address 0x05d0
		x"1af6", x"0225", x"0037", x"c285", x"050a", x"06a0", x"061c", x"3700", -- address 0x05e0
		x"04c5", x"2fa0", x"0128", x"8040", x"1304", x"04c3", x"2fa0", x"0137", -- address 0x05f0
		x"10e2", x"2fa0", x"012b", x"0203", x"003c", x"2fa0", x"0134", x"0603", -- address 0x0600
		x"16fc", x"0720", x"ec46", x"2fa0", x"00f2", x"104a", x"c13b", x"2f04", -- address 0x0610
		x"0984", x"a144", x"2e8a", x"0223", x"0005", x"0204", x"0004", x"0b4a", -- address 0x0620
		x"c30a", x"09cc", x"a14c", x"0225", x"0030", x"028c", x"000a", x"1a02", -- address 0x0630
		x"0225", x"0007", x"0604", x"16f3", x"045b", x"2fa0", x"002d", x"2f44", -- address 0x0640
		x"0284", x"5900", x"162d", x"0206", x"1100", x"2f06", x"04c7", x"04c8", -- address 0x0650
		x"06a0", x"0728", x"100b", x"d22a", x"070e", x"132d", x"06a0", x"0722", -- address 0x0660
		x"100e", x"0205", x"0008", x"0878", x"0468", x"0678", x"0286", x"0047", -- address 0x0670
		x"1106", x"0286", x"004a", x"1516", x"0226", x"ffc9", x"10ec", x"0286", -- address 0x0680
		x"003a", x"1610", x"04ca", x"0705", x"020c", x"0080", x"1f0f", x"16fb", -- address 0x0690
		x"0605", x"16fc", x"c28a", x"1609", x"2fa0", x"00f2", x"2fa0", x"ec02", -- address 0x06a0
		x"0460", x"0142", x"04c0", x"070a", x"10ee", x"c000", x"1302", x"0460", -- address 0x06b0
		x"0208", x"0460", x"0204", x"2f46", x"9806", x"00f2", x"16fc", x"10c6", -- address 0x06c0
		x"a280", x"c24a", x"10c4", x"a280", x"ce4a", x"10c1", x"a1ca", x"13bf", -- address 0x06d0
		x"0200", x"0001", x"10e8", x"020a", x"ec02", x"1003", x"0645", x"020a", -- address 0x06e0
		x"ec22", x"2f46", x"de86", x"0986", x"a1c6", x"0605", x"16fa", x"10af", -- address 0x06f0
		x"a280", x"c38a", x"10ac", x"024a", x"fffe", x"c00a", x"10a8", x"3745", -- address 0x0700
		x"443a", x"3a3a", x"3a32", x"f22d", x"2c30", x"2f47", x"1e00", x"3a3a", -- address 0x0710
		x"3bf3", x"0205", x"fffc", x"1001", x"0705", x"04ca", x"2f46", x"0286", -- address 0x0720
		x"2000", x"11fc", x"0286", x"5f00", x"15f9", x"0986", x"0288", x"3200", -- address 0x0730
		x"1301", x"a1c6", x"0286", x"0030", x"1112", x"0286", x"0039", x"1208", -- address 0x0740
		x"0286", x"0041", x"110c", x"0286", x"0046", x"1509", x"0226", x"0009", -- address 0x0750
		x"0246", x"000f", x"0a4a", x"a286", x"0585", x"16e0", x"05cb", x"045b", -- address 0x0760
		x"0203", x"8402", x"0204", x"05c0", x"0a25", x"1103", x"4008", x"4048", -- address 0x0770
		x"1007", x"0223", x"1000", x"0224", x"ffc0", x"0a82", x"1001", x"0484", -- address 0x0780
		x"0483", x"1603", x"2fa0", x"00f2", x"2e80", x"8040", x"16f8", x"0459", -- address 0x0790
		x"2fa0", x"00c0", x"c100", x"a101", x"2e84", x"2fa0", x"00c9", x"6001", -- address 0x07a0
		x"2e80", x"0459", x"0560", x"ec44", x"0459", x"04e0", x"ec4e", x"04e0", -- address 0x07b0
		x"ec4c", x"c240", x"2fa0", x"00f2", x"020a", x"0850", x"0200", x"ec52", -- address 0x07c0
		x"0208", x"0006", x"04f0", x"0608", x"15fd", x"2e89", x"2fa0", x"001c", -- address 0x07d0
		x"069a", x"0284", x"0020", x"1316", x"0284", x"002a", x"1605", x"069a", -- address 0x07e0
		x"0284", x"000d", x"16fc", x"10e6", x"06a0", x"0bee", x"c807", x"ec52", -- address 0x07f0
		x"c809", x"ec54", x"c107", x"06a0", x"0c64", x"1321", x"9807", x"0bf3", -- address 0x0800
		x"1303", x"1004", x"2fa0", x"0021", x"2fa0", x"0021", x"0207", x"0ce3", -- address 0x0810
		x"04c5", x"04c6", x"069a", x"06a0", x"0c34", x"1643", x"0ab4", x"0587", -- address 0x0820
		x"d017", x"1102", x"1372", x"05c6", x"0a10", x"09e0", x"8005", x"11f7", -- address 0x0830
		x"156c", x"d017", x"0a30", x"9100", x"16f2", x"0585", x"10eb", x"1065", -- address 0x0840
		x"2f44", x"0284", x"1b00", x"13b6", x"0284", x"2000", x"1a01", x"2f04", -- address 0x0850
		x"0984", x"c804", x"ec60", x"045b", x"069a", x"0284", x"0027", x"1655", -- address 0x0860
		x"c1c9", x"75d7", x"0588", x"069a", x"0284", x"0027", x"1358", x"06c4", -- address 0x0870
		x"ddc4", x"10f7", x"06a0", x"0b14", x"c806", x"ec54", x"1064", x"070e", -- address 0x0880
		x"c006", x"06a0", x"0b14", x"c809", x"ec54", x"0280", x"0014", x"1605", -- address 0x0890
		x"a189", x"1303", x"0586", x"8246", x"1a38", x"c246", x"0249", x"fffe", -- address 0x08a0
		x"1052", x"c145", x"13af", x"d017", x"1130", x"070e", x"0286", x"0032", -- address 0x08b0
		x"13e1", x"0286", x"009a", x"13d0", x"c026", x"0d76", x"c040", x"0241", -- address 0x08c0
		x"fff0", x"1302", x"c641", x"05c8", x"c040", x"0241", x"000f", x"d021", -- address 0x08d0
		x"0cd6", x"06c0", x"0260", x"ffe0", x"c040", x"0921", x"0241", x"0006", -- address 0x08e0
		x"c061", x"0cc6", x"1307", x"0284", x"0020", x"160f", x"04ce", x"020f", -- address 0x08f0
		x"0904", x"0691", x"c040", x"0ad1", x"09c1", x"c061", x"0cc6", x"1309", -- address 0x0900
		x"04c0", x"04ce", x"020f", x"0922", x"0691", x"2fa0", x"00d1", x"0460", -- address 0x0910
		x"07c4", x"0284", x"000d", x"1307", x"0284", x"0020", x"16f6", x"069a", -- address 0x0920
		x"0284", x"000d", x"16fc", x"0280", x"0030", x"135c", x"2f20", x"00f2", -- address 0x0930
		x"2e89", x"c089", x"06a0", x"0c86", x"0204", x"2052", x"c0c3", x"1301", -- address 0x0940
		x"06c4", x"2f04", x"2eb9", x"2fa0", x"00f2", x"0648", x"15f1", x"0200", -- address 0x0950
		x"ec56", x"06a0", x"0c9a", x"06a0", x"0c9a", x"c120", x"ec52", x"1331", -- address 0x0960
		x"0224", x"8000", x"06a0", x"0c64", x"1608", x"06a0", x"09d6", x"c390", -- address 0x0970
		x"c403", x"06a0", x"09e6", x"c00e", x"16fa", x"0224", x"8080", x"06a0", -- address 0x0980
		x"0c64", x"161a", x"06a0", x"09d6", x"04ce", x"0580", x"d390", x"c083", -- address 0x0990
		x"6080", x"0602", x"0a72", x"1907", x"0600", x"2e80", x"2fa0", x"00d1", -- address 0x09a0
		x"2fa0", x"00f2", x"1004", x"d402", x"0600", x"06a0", x"09e6", x"087e", -- address 0x09b0
		x"05ce", x"1302", x"a00e", x"10e8", x"0200", x"ec52", x"04c4", x"06a0", -- address 0x09c0
		x"0c9c", x"0460", x"07c8", x"c012", x"04e2", x"fffe", x"0620", x"ec4c", -- address 0x09d0
		x"c0e0", x"ec54", x"045b", x"2e80", x"2f20", x"0a05", x"2e90", x"2fa0", -- address 0x09e0
		x"00f2", x"045b", x"2fa0", x"001f", x"2ea0", x"ec4c", x"0460", x"0142", -- address 0x09f0
		x"069a", x"0284", x"002a", x"131a", x"0284", x"0040", x"1622", x"06a0", -- address 0x0a00
		x"0b14", x"c088", x"a089", x"c486", x"05c8", x"0206", x"0020", x"0284", -- address 0x0a10
		x"0028", x"1608", x"06a0", x"0ad0", x"0266", x"0020", x"0284", x"0029", -- address 0x0a20
		x"1649", x"069a", x"c000", x"1601", x"0a66", x"1040", x"06a0", x"0ad0", -- address 0x0a30
		x"0266", x"0010", x"0284", x"002b", x"1603", x"069a", x"0266", x"0030", -- address 0x0a40
		x"10f1", x"020e", x"0a34", x"c80e", x"ec5e", x"0460", x"0ad6", x"06a0", -- address 0x0a50
		x"0ad0", x"0a46", x"102b", x"c006", x"0280", x"0030", x"1604", x"0284", -- address 0x0a60
		x"000d", x"1312", x"070e", x"06a0", x"0b14", x"0280", x"0030", x"130b", -- address 0x0a70
		x"c089", x"a088", x"c486", x"05c8", x"0280", x"0026", x"1605", x"070e", -- address 0x0a80
		x"0284", x"002c", x"13f0", x"c386", x"045f", x"06a0", x"0ad0", x"10ca", -- address 0x0a90
		x"06a0", x"0b14", x"c089", x"05c2", x"6182", x"0816", x"0286", x"007f", -- address 0x0aa0
		x"1507", x"0286", x"ff80", x"1104", x"0246", x"00ff", x"e646", x"045f", -- address 0x0ab0
		x"2fa0", x"00d6", x"0460", x"091a", x"070e", x"06a0", x"0b14", x"10ee", -- address 0x0ac0
		x"c80b", x"ec5e", x"069a", x"020c", x"0b04", x"0284", x"0052", x"130c", -- address 0x0ad0
		x"0284", x"003a", x"110a", x"0284", x"003e", x"1309", x"020e", x"fffe", -- address 0x0ae0
		x"020d", x"0b04", x"0460", x"0b18", x"069a", x"0460", x"0c2a", x"069a", -- address 0x0af0
		x"0460", x"0c0c", x"c145", x"11de", x"0286", x"0010", x"14db", x"c2e0", -- address 0x0b00
		x"ec5e", x"045b", x"c34b", x"069a", x"04e0", x"ec50", x"0284", x"0027", -- address 0x0b10
		x"1307", x"0284", x"002d", x"1610", x"054d", x"05ce", x"069a", x"1011", -- address 0x0b20
		x"04c6", x"04ce", x"069a", x"0284", x"0027", x"1304", x"06c6", x"d106", -- address 0x0b30
		x"c184", x"10f8", x"069a", x"1043", x"0284", x"002b", x"13ee", x"c38e", -- address 0x0b40
		x"154b", x"0284", x"0024", x"1603", x"c189", x"069a", x"1037", x"0284", -- address 0x0b50
		x"003e", x"1604", x"069a", x"06a0", x"0c0a", x"1030", x"06a0", x"0c34", -- address 0x0b60
		x"11a9", x"1325", x"06a0", x"0c28", x"1029", x"c38e", x"16a3", x"c059", -- address 0x0b70
		x"04c2", x"06a0", x"0c86", x"c4c9", x"0241", x"f000", x"0281", x"1000", -- address 0x0b80
		x"1611", x"0264", x"0080", x"c189", x"0643", x"c4c4", x"8820", x"ec56", -- address 0x0b90
		x"ec5a", x"1603", x"c1a0", x"ec58", x"1012", x"06a0", x"0c64", x"1601", -- address 0x0ba0
		x"c192", x"100d", x"a4c8", x"0264", x"8000", x"04c6", x"10ed", x"06a0", -- address 0x0bb0
		x"0bee", x"c107", x"06a0", x"0c64", x"16d8", x"c192", x"05ce", x"c120", -- address 0x0bc0
		x"ec60", x"c34d", x"1502", x"0506", x"054d", x"c145", x"1194", x"c38e", -- address 0x0bd0
		x"1305", x"a806", x"ec50", x"109d", x"c1a0", x"ec50", x"045d", x"c30b", -- address 0x0be0
		x"0207", x"0031", x"06a0", x"0c34", x"111c", x"1303", x"0a87", x"1919", -- address 0x0bf0
		x"1001", x"0a87", x"a1c4", x"069a", x"10f5", x"c30b", x"0202", x"0010", -- address 0x0c00
		x"04c6", x"0705", x"06a0", x"0c34", x"110c", x"8083", x"1409", x"c146", -- address 0x0c10
		x"3942", x"a183", x"069a", x"10f6", x"c30b", x"0202", x"000a", x"10f0", -- address 0x0c20
		x"0705", x"045c", x"0701", x"c0c4", x"0284", x"0024", x"1306", x"0223", -- address 0x0c30
		x"ffd0", x"170e", x"0283", x"0009", x"1502", x"0501", x"045b", x"0223", -- address 0x0c40
		x"fff9", x"0283", x"000a", x"1a04", x"0283", x"0023", x"1b01", x"04c1", -- address 0x0c50
		x"c041", x"045b", x"0703", x"c060", x"ec4e", x"130b", x"0a21", x"0202", -- address 0x0c60
		x"ec62", x"a042", x"04c3", x"05c2", x"8c84", x"1303", x"8042", x"1afb", -- address 0x0c70
		x"0583", x"c0c3", x"045b", x"0203", x"ec58", x"84c2", x"1305", x"0203", -- address 0x0c80
		x"ec5c", x"84c2", x"1301", x"04c3", x"045b", x"c110", x"c30b", x"06a0", -- address 0x0c90
		x"0c64", x"130d", x"c104", x"1304", x"04c4", x"05a0", x"ec4c", x"10f7", -- address 0x0ca0
		x"05a0", x"ec4e", x"c0a0", x"ec4e", x"0a22", x"0222", x"ec62", x"0642", -- address 0x0cb0
		x"ccb0", x"c4b0", x"045c", x"0000", x"0a00", x"0a9a", x"0a66", x"0a5e", -- address 0x0cc0
		x"0aa0", x"0ac8", x"088e", x"0905", x"0a0a", x"1408", x"0013", x"0a06", -- address 0x0cd0
		x"0310", x"0307", x"0122", x"5329", x"aec4", x"69af", x"d267", x"022c", -- address 0x0ce0
		x"d770", x"b353", x"0322", x"29ab", x"cf6e", x"66ac", x"52af", x"43ba", -- address 0x0cf0
		x"4384", x"a1d4", x"61a5", x"4374", x"a956", x"7385", x"ae44", x"b155", -- address 0x0d00
		x"89a4", x"cc65", x"ae43", x"7456", x"8aa5", x"51a7", x"5428", x"452c", -- address 0x0d10
		x"4554", x"ad50", x"ae43", x"454f", x"af43", x"508c", x"a4c3", x"7229", -- address 0x0d20
		x"cd69", x"b2c5", x"78b3", x"54b7", x"5069", x"8daf", x"5662", x"b059", -- address 0x0d30
		x"738e", x"a547", x"af50", x"8fb2", x"4992", x"b3c5", x"74b4", x"d770", -- address 0x0d40
		x"1322", x"4f5a", x"a5d4", x"6fac", x"41af", x"4362", x"b241", x"434c", -- address 0x0d50
		x"b4c3", x"72d3", x"74d7", x"70b7", x"d062", x"ba43", x"6294", x"22a5", -- address 0x0d60
		x"d874", x"18af", x"5052", x"0000", x"a000", x"b000", x"0745", x"0227", -- address 0x0d70
		x"0247", x"000d", x"0445", x"0685", x"0405", x"000d", x"8000", x"9000", -- address 0x0d80
		x"0287", x"03a6", x"03c6", x"04c5", x"2002", x"2402", x"000a", x"0605", -- address 0x0d90
		x"0645", x"3c08", x"0185", x"000c", x"0006", x"0346", x"0585", x"05c5", -- address 0x0da0
		x"0545", x"1301", x"1501", x"1b01", x"1401", x"1a01", x"1201", x"1101", -- address 0x0db0
		x"1001", x"1701", x"1601", x"1901", x"1801", x"1c01", x"3003", x"0207", -- address 0x0dc0
		x"030a", x"03e6", x"008b", x"009b", x"02ea", x"c000", x"d000", x"3808", -- address 0x0dd0
		x"01c5", x"0505", x"1006", x"0267", x"0366", x"0386", x"6000", x"7000", -- address 0x0de0
		x"1d09", x"1e09", x"0705", x"0a04", x"e000", x"f000", x"0804", x"0b04", -- address 0x0df0
		x"0904", x"3403", x"02cb", x"02ab", x"06c5", x"4000", x"5000", x"1f09", -- address 0x0e00
		x"0006", x"0485", x"2c08", x"2802", x"0000", x"02e0", x"ec00", x"0203", -- address 0x0e10
		x"ec4c", x"0205", x"ed00", x"0206", x"effe", x"ccc5", x"ccc6", x"ccc5", -- address 0x0e20
		x"04c5", x"04d3", x"0209", x"ec2e", x"c820", x"ec44", x"ec54", x"020c", -- address 0x0e30
		x"0400", x"1d1f", x"3220", x"013b", x"1e0d", x"3320", x"0096", x"1d10", -- address 0x0e40
		x"020c", x"0000", x"1d0e", x"3220", x"013b", x"04c1", x"04c2", x"c660", -- address 0x0e50
		x"013e", x"2fa0", x"00e3", x"05e0", x"ec44", x"020c", x"0000", x"1f15", -- address 0x0e60
		x"1334", x"020c", x"0400", x"1f15", x"1303", x"c041", x"162c", x"10f5", -- address 0x0e70
		x"c660", x"0140", x"c082", x"1625", x"2f4a", x"028a", x"0000", x"13ed", -- address 0x0e80
		x"028a", x"7f00", x"13ea", x"028a", x"1000", x"160d", x"2f4a", x"028a", -- address 0x0e90
		x"0000", x"13fc", x"028a", x"3700", x"130e", x"028a", x"3c00", x"16dd", -- address 0x0ea0
		x"2f20", x"013c", x"10da", x"028a", x"1200", x"1602", x"0460", x"1070", -- address 0x0eb0
		x"028a", x"1100", x"1602", x"0460", x"0fa0", x"c660", x"013e", x"2f0a", -- address 0x0ec0
		x"10cc", x"0460", x"107c", x"0460", x"0fc8", x"c660", x"013e", x"2f4a", -- address 0x0ed0
		x"028a", x"1a00", x"1605", x"c820", x"ec54", x"ec44", x"0460", x"0142", -- address 0x0ee0
		x"028a", x"0300", x"1310", x"028a", x"1200", x"13e0", x"028a", x"1400", -- address 0x0ef0
		x"1602", x"0460", x"10fe", x"c041", x"16e6", x"c082", x"16e2", x"c660", -- address 0x0f00
		x"0140", x"2f0a", x"10aa", x"c660", x"013e", x"c820", x"ec54", x"ec44", -- address 0x0f10
		x"2fa0", x"00d8", x"2eca", x"2fa0", x"00de", x"06a0", x"0f42", x"5500", -- address 0x0f20
		x"0f7e", x"4400", x"0f94", x"5400", x"0f5a", x"5100", x"0e5a", x"0000", -- address 0x0f30
		x"05cb", x"c01b", x"1304", x"82bb", x"16fb", x"c2db", x"045b", x"2fa0", -- address 0x0f40
		x"00f5", x"10e1", x"2fa0", x"00ff", x"10de", x"2e4a", x"0f16", x"0f54", -- address 0x0f50
		x"0a2a", x"064a", x"12f7", x"028a", x"0023", x"14f4", x"020c", x"0400", -- address 0x0f60
		x"1d0b", x"1d0c", x"332a", x"0084", x"1e0b", x"1e0c", x"10cc", x"2e4a", -- address 0x0f70
		x"0f88", x"0f54", x"c80a", x"ec50", x"2e4a", x"0f16", x"0f54", x"c80a", -- address 0x0f80
		x"ec4e", x"10c1", x"2e4a", x"0f16", x"0f54", x"c80a", x"ec4c", x"10bb", -- address 0x0f90
		x"0701", x"c1e0", x"ec52", x"112d", x"1533", x"c1e0", x"ec50", x"8807", -- address 0x0fa0
		x"ec4e", x"1b37", x"c660", x"0140", x"04c5", x"04c3", x"2fa0", x"0137", -- address 0x0fb0
		x"c287", x"06a0", x"1042", x"3900", x"c297", x"06a0", x"1042", x"4200", -- address 0x0fc0
		x"8807", x"ec4e", x"1a03", x"0720", x"ec52", x"1004", x"05c7", x"0283", -- address 0x0fd0
		x"003c", x"111d", x"0225", x"0037", x"c285", x"050a", x"06a0", x"1042", -- address 0x0fe0
		x"3700", x"c807", x"ec50", x"2fa0", x"0128", x"c160", x"ec54", x"110e", -- address 0x0ff0
		x"10cf", x"2fa0", x"0137", x"2fa0", x"00e0", x"05e0", x"ec52", x"10f5", -- address 0x1000
		x"2fa0", x"0137", x"2fa0", x"0131", x"04e0", x"ec52", x"04c1", x"0460", -- address 0x1010
		x"0e6a", x"2fa0", x"0137", x"2fa0", x"0131", x"c660", x"013e", x"c820", -- address 0x1020
		x"ec54", x"ec44", x"2fa0", x"011f", x"05e0", x"ec44", x"0720", x"ec4c", -- address 0x1030
		x"10eb", x"c03b", x"2f00", x"0980", x"a140", x"2e8a", x"0223", x"0005", -- address 0x1040
		x"0200", x"0004", x"0b4a", x"c18a", x"09c6", x"a146", x"0225", x"0030", -- address 0x1050
		x"0286", x"000a", x"1a02", x"0225", x"0007", x"0600", x"16f3", x"045b", -- address 0x1060
		x"0702", x"c660", x"0140", x"c020", x"ec4c", x"04c7", x"2f46", x"0286", -- address 0x1070
		x"1400", x"133d", x"c220", x"ec52", x"1657", x"0286", x"2000", x"11f6", -- address 0x1080
		x"0286", x"5f00", x"15f3", x"0705", x"04ca", x"06a0", x"073a", x"100b", -- address 0x1090
		x"d22a", x"1152", x"1332", x"06a0", x"0722", x"100e", x"0205", x"0008", -- address 0x10a0
		x"0878", x"0468", x"10b2", x"0286", x"0047", x"1106", x"0286", x"004a", -- address 0x10b0
		x"1522", x"0226", x"ffc9", x"10ec", x"0286", x"003a", x"161c", x"103e", -- address 0x10c0
		x"020c", x"0400", x"04c5", x"1f0f", x"16fd", x"0605", x"16fc", x"c660", -- address 0x10d0
		x"013e", x"c820", x"ec54", x"ec44", x"0720", x"ec4c", x"c000", x"1303", -- address 0x10e0
		x"2fa0", x"010a", x"1002", x"2fa0", x"0115", x"05e0", x"ec44", x"04c2", -- address 0x10f0
		x"04e0", x"ec52", x"1021", x"04c0", x"10e3", x"2f46", x"9806", x"00f2", -- address 0x1100
		x"16fc", x"04c7", x"1019", x"a1ca", x"1317", x"0700", x"10d9", x"a280", -- address 0x1110
		x"c0ca", x"1012", x"a280", x"ccca", x"100f", x"0645", x"2f46", x"0986", -- address 0x1120
		x"13fd", x"a1c6", x"0605", x"16fa", x"1007", x"a280", x"c80a", x"ec1c", -- address 0x1130
		x"1003", x"024a", x"fffe", x"c00a", x"0460", x"0e6a", x"0720", x"ec52", -- address 0x1140
		x"10fb", x"3d45", x"443c", x"3c3c", x"3c32", x"e437", x"363a", x"3948", -- address 0x1150
		x"2a00", x"3c3c", x"3d8b", x"c141", x"0208", x"12d8", x"0209", x"12ba", -- address 0x1160
		x"0207", x"12a6", x"2fa0", x"00f2", x"0206", x"202c", x"c050", x"2e80", -- address 0x1170
		x"2f06", x"2e81", x"2f06", x"04c3", x"c050", x"0241", x"fff0", x"c2a3", -- address 0x1180
		x"13b4", x"c08a", x"1329", x"024a", x"fff0", x"8281", x"1402", x"0643", -- address 0x1190
		x"10f6", x"c050", x"0a13", x"0223", x"14d6", x"604a", x"0242", x"000f", -- address 0x11a0
		x"d0a2", x"11ba", x"0972", x"0462", x"11ba", x"060c", x"061f", x"232b", -- address 0x11b0
		x"3337", x"063f", x"4145", x"0697", x"0698", x"2f06", x"0961", x"0698", -- address 0x11c0
		x"103d", x"c041", x"1603", x"0203", x"14da", x"1024", x"06c1", x"0871", -- address 0x11d0
		x"05c1", x"a040", x"0697", x"1004", x"c050", x"0203", x"14de", x"0697", -- address 0x11e0
		x"2f20", x"14f5", x"2e81", x"102a", x"0697", x"0698", x"c209", x"10e5", -- address 0x11f0
		x"d041", x"16f2", x"0b41", x"d081", x"0a61", x"09c2", x"a042", x"10f4", -- address 0x1200
		x"8810", x"1320", x"1603", x"0203", x"14ee", x"1004", x"0697", x"10d7", -- address 0x1210
		x"c041", x"16e2", x"0697", x"1012", x"0ac1", x"18de", x"09c1", x"0697", -- address 0x1220
		x"0698", x"2f06", x"c070", x"10dc", x"0697", x"1019", x"c041", x"16d4", -- address 0x1230
		x"0697", x"10f8", x"0ac1", x"18d0", x"09c1", x"10e2", x"c145", x"1603", -- address 0x1240
		x"c740", x"0460", x"0142", x"c320", x"013e", x"1f15", x"1604", x"2f42", -- address 0x1250
		x"0282", x"2f00", x"13f5", x"8140", x"1bf3", x"0460", x"1168", x"0203", -- address 0x1260
		x"2d31", x"06c1", x"0881", x"1315", x"1502", x"2f03", x"0501", x"0281", -- address 0x1270
		x"0064", x"1104", x"0a83", x"2f03", x"0221", x"ff9c", x"0204", x"000a", -- address 0x1280
		x"c081", x"04c1", x"3c44", x"0a83", x"1302", x"c041", x"1301", x"0699", -- address 0x1290
		x"c042", x"0699", x"10d3", x"0202", x"0004", x"2f13", x"0583", x"0602", -- address 0x12a0
		x"16fc", x"2f06", x"06c6", x"05c0", x"045b", x"c0c1", x"0ac3", x"0943", -- address 0x12b0
		x"0283", x"0900", x"1203", x"06c3", x"0223", x"0126", x"0223", x"3000", -- address 0x12c0
		x"2f03", x"0a83", x"16fd", x"045b", x"0204", x"2a52", x"c081", x"0aa2", -- address 0x12d0
		x"09e2", x"1603", x"06c4", x"2f04", x"10e8", x"0602", x"1602", x"2f04", -- address 0x12e0
		x"10f9", x"0602", x"1610", x"2fa0", x"14f4", x"2eb0", x"c081", x"0ac2", -- address 0x12f0
		x"13ea", x"0202", x"2829", x"2f02", x"06c4", x"2f04", x"c30b", x"0699", -- address 0x1300
		x"06c2", x"2f02", x"045c", x"2fa0", x"14f7", x"0202", x"002b", x"10f6", -- address 0x1310
		x"045b", x"0000", x"008b", x"009b", x"0185", x"01c5", x"0207", x"0227", -- address 0x1320
		x"0247", x"0267", x"0287", x"02ab", x"02cb", x"02ea", x"030a", x"0346", -- address 0x1330
		x"0366", x"0386", x"03a6", x"03c6", x"03e6", x"0405", x"0445", x"0485", -- address 0x1340
		x"04c5", x"0505", x"0545", x"0585", x"05c5", x"0605", x"0645", x"0685", -- address 0x1350
		x"06c5", x"0705", x"0745", x"0804", x"0904", x"0a04", x"0b04", x"1001", -- address 0x1360
		x"1101", x"1201", x"1301", x"1401", x"1501", x"1601", x"1701", x"1801", -- address 0x1370
		x"1901", x"1a01", x"1b01", x"1c01", x"1d09", x"1e09", x"1f09", x"2002", -- address 0x1380
		x"2402", x"2802", x"2c03", x"3003", x"3403", x"3808", x"3c08", x"4000", -- address 0x1390
		x"5000", x"6000", x"7000", x"8000", x"9000", x"a000", x"b000", x"c000", -- address 0x13a0
		x"d000", x"e000", x"f000", x"4c53", x"5420", x"4c57", x"5020", x"4449", -- address 0x13b0
		x"5653", x"4d50", x"5953", x"4c49", x"2020", x"4149", x"2020", x"414e", -- address 0x13c0
		x"4449", x"4f52", x"4920", x"4349", x"2020", x"5354", x"5750", x"5354", -- address 0x13d0
		x"5354", x"4c57", x"5049", x"4c49", x"4d49", x"4944", x"4c45", x"5253", -- address 0x13e0
		x"4554", x"5254", x"5750", x"434b", x"4f4e", x"434b", x"4f46", x"4c52", -- address 0x13f0
		x"4558", x"424c", x"5750", x"4220", x"2020", x"5820", x"2020", x"434c", -- address 0x1400
		x"5220", x"4e45", x"4720", x"494e", x"5620", x"494e", x"4320", x"494e", -- address 0x1410
		x"4354", x"4445", x"4320", x"4445", x"4354", x"424c", x"2020", x"5357", -- address 0x1420
		x"5042", x"5345", x"544f", x"4142", x"5320", x"5352", x"4120", x"5352", -- address 0x1430
		x"4c20", x"534c", x"4120", x"5352", x"4320", x"4a4d", x"5020", x"4a4c", -- address 0x1440
		x"5420", x"4a4c", x"4520", x"4a45", x"5120", x"4a48", x"4520", x"4a47", -- address 0x1450
		x"5420", x"4a4e", x"4520", x"4a4e", x"4320", x"4a4f", x"4320", x"4a4e", -- address 0x1460
		x"4f20", x"4a4c", x"2020", x"4a48", x"2020", x"4a4f", x"5020", x"5342", -- address 0x1470
		x"4f20", x"5342", x"5a20", x"5442", x"2020", x"434f", x"4320", x"435a", -- address 0x1480
		x"4320", x"584f", x"5220", x"584f", x"5020", x"4c44", x"4352", x"5354", -- address 0x1490
		x"4352", x"4d50", x"5920", x"4449", x"5620", x"535a", x"4320", x"535a", -- address 0x14a0
		x"4342", x"5320", x"2020", x"5342", x"2020", x"4320", x"2020", x"4342", -- address 0x14b0
		x"2020", x"4120", x"2020", x"4142", x"2020", x"4d4f", x"5620", x"4d4f", -- address 0x14c0
		x"5642", x"534f", x"4320", x"534f", x"4342", x"4e4f", x"5020", x"4441", -- address 0x14d0
		x"5441", x"5445", x"5854", x"414f", x"5247", x"454e", x"4420", x"5254", -- address 0x14e0
		x"2020", x"0000", x"403e", x"002a", x"5200", x"ffff", x"ffff", x"ffff", -- address 0x14f0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1500
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1510
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1520
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1530
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1540
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1550
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1560
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1570
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1580
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1590
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x15a0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x15b0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x15c0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x15d0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x15e0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x15f0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1600
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1610
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1620
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1630
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1640
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1650
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1660
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1670
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1680
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1690
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x16a0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x16b0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x16c0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x16d0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x16e0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x16f0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1700
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1710
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1720
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1730
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1740
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1750
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1760
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1770
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1780
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1790
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x17a0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x17b0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x17c0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x17d0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x17e0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x17f0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1800
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1810
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1820
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1830
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1840
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1850
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1860
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1870
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1880
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1890
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x18a0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x18b0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x18c0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x18d0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x18e0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x18f0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1900
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1910
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1920
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1930
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1940
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1950
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1960
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1970
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1980
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1990
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x19a0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x19b0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x19c0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x19d0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x19e0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x19f0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1a00
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1a10
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1a20
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1a30
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1a40
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1a50
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1a60
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1a70
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1a80
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1a90
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1aa0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1ab0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1ac0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1ad0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1ae0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1af0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1b00
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1b10
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1b20
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1b30
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1b40
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1b50
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1b60
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1b70
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1b80
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1b90
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1ba0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1bb0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1bc0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1bd0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1be0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1bf0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1c00
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1c10
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1c20
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1c30
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1c40
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1c50
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1c60
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1c70
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1c80
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1c90
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1ca0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1cb0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1cc0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1cd0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1ce0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1cf0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1d00
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1d10
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1d20
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1d30
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1d40
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1d50
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1d60
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1d70
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1d80
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1d90
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1da0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1db0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1dc0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1dd0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1de0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1df0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1e00
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1e10
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1e20
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1e30
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1e40
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1e50
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1e60
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1e70
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1e80
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1e90
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1ea0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1eb0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1ec0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1ed0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1ee0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1ef0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1f00
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1f10
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1f20
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1f30
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1f40
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1f50
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1f60
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1f70
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1f80
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1f90
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1fa0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1fb0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1fc0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1fd0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", -- address 0x1fe0
		x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff"  -- address 0x1ff0
   );

begin

	process(CLK, nCS)
	variable idx : integer range 0 to size;
	begin
		if rising_edge(CLK) and nCS='0' then
			idx := to_integer( unsigned( ADDR ));
			DO <= rom( idx );
		end if;
	end process;

end rom_arch;

