----------------------------------------------------------------------------------
-- Engineer:	Erik Piehl 
-- 
-- Create Date:    07:01:30 04/15/2017 
-- Design Name: 	 testrom.vhd
-- Module Name:    testrom - Behavioral 
-- Project Name: 	 TMS9900 Test ROM code
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity testrom is
    Port ( clk : in  STD_LOGIC;
           addr : in  STD_LOGIC_VECTOR (11 downto 0);
           data_out : out  STD_LOGIC_VECTOR (15 downto 0));
end testrom;

architecture Behavioral of testrom is
	constant romLast : integer := 16383;
	type pgmRomArray is array(0 to romLast) of STD_LOGIC_VECTOR (15 downto 0);
	constant pgmRom : pgmRomArray := (  
            x"ec00"
           ,x"0226" -- 0002
           ,x"f0d6" -- 0004
           ,x"f0f6" -- 0006
           ,x"f0ca" -- 0008
           ,x"f0ea" -- 000A
           ,x"f0be" -- 000C
           ,x"f0de" -- 000E
           ,x"f0b2" -- 0010
           ,x"f0d2" -- 0012
           ,x"0d0a" -- 0014
           ,x"4d4f" -- 0016
           ,x"4e3f" -- 0018
           ,x"2000" -- 001A
           ,x"2020" -- 001C
           ,x"2020" -- 001E
           ,x"2020" -- 0020
           ,x"000d" -- 0022
           ,x"0a42" -- 0024
           ,x"5000" -- 0026
           ,x"4944" -- 0028
           ,x"543d" -- 002A
           ,x"000d" -- 002C
           ,x"0a52" -- 002E
           ,x"4541" -- 0030
           ,x"4459" -- 0032
           ,x"2059" -- 0034
           ,x"2f4e" -- 0036
           ,x"2000" -- 0038
           ,x"5700" -- 003A
           ,x"5000" -- 003C
           ,x"5300" -- 003E
           ,x"f0ac" -- 0040
           ,x"f0be" -- 0042
           ,x"f09e" -- 0044
           ,x"f0b0" -- 0046
           ,x"f090" -- 0048
           ,x"f0a2" -- 004A
           ,x"f082" -- 004C
           ,x"f094" -- 004E
           ,x"f074" -- 0050
           ,x"f086" -- 0052
           ,x"f066" -- 0054
           ,x"f078" -- 0056
           ,x"f058" -- 0058
           ,x"f06a" -- 005A
           ,x"f04a" -- 005C
           ,x"f05c" -- 005E
           ,x"ec24" -- 0060
           ,x"03f8" -- 0062
           ,x"ec24" -- 0064
           ,x"0396" -- 0066
           ,x"ec24" -- 0068
           ,x"0402" -- 006A
           ,x"ec0a" -- 006C
           ,x"0326" -- 006E
           ,x"ec16" -- 0070
           ,x"02ee" -- 0072
           ,x"ec16" -- 0074
           ,x"02e2" -- 0076
           ,x"ec24" -- 0078
           ,x"032c" -- 007A
           ,x"ec00" -- 007C
           ,x"0442" -- 007E
           ,x"0460" -- 0080
           ,x"0142" -- 0082
           ,x"0009" -- 0084
           ,x"001a" -- 0086
           ,x"0012" -- 0088
           ,x"0034" -- 008A
           ,x"0023" -- 008C
           ,x"0068" -- 008E
           ,x"0046" -- 0090
           ,x"00d0" -- 0092
           ,x"008d" -- 0094
           ,x"01a1" -- 0096
           ,x"0119" -- 0098
           ,x"0341" -- 009A
           ,x"02a4" -- 009C
           ,x"04d0" -- 009E
           ,x"7fff" -- 00A0
           ,x"0638" -- 00A2
           ,x"0d0a" -- 00A4
           ,x"4552" -- 00A6
           ,x"524f" -- 00A8
           ,x"5220" -- 00AA
           ,x"000d" -- 00AC
           ,x"0a45" -- 00AE
           ,x"564d" -- 00B0
           ,x"4255" -- 00B2
           ,x"4720" -- 00B4
           ,x"2052" -- 00B6
           ,x"312e" -- 00B8
           ,x"3000" -- 00BA
           ,x"0d0a" -- 00BC
           ,x"5200" -- 00BE
           ,x"0d0a" -- 00C0
           ,x"4831" -- 00C2
           ,x"2b48" -- 00C4
           ,x"323d" -- 00C6
           ,x"0020" -- 00C8
           ,x"4831" -- 00CA
           ,x"2d48" -- 00CC
           ,x"323d" -- 00CE
           ,x"0020" -- 00D0
           ,x"4552" -- 00D2
           ,x"524f" -- 00D4
           ,x"5200" -- 00D6
           ,x"0d0a" -- 00D8
           ,x"434f" -- 00DA
           ,x"4d3f" -- 00DC
           ,x"2000" -- 00DE
           ,x"3a0d" -- 00E0
           ,x"000d" -- 00E2
           ,x"0a54" -- 00E4
           ,x"4552" -- 00E6
           ,x"4d49" -- 00E8
           ,x"4e41" -- 00EA
           ,x"4c20" -- 00EC
           ,x"4d4f" -- 00EE
           ,x"4445" -- 00F0
           ,x"0d0a" -- 00F2
           ,x"000d" -- 00F4
           ,x"0a43" -- 00F6
           ,x"4d44" -- 00F8
           ,x"2045" -- 00FA
           ,x"5252" -- 00FC
           ,x"000d" -- 00FE
           ,x"0a50" -- 0100
           ,x"4152" -- 0102
           ,x"4d20" -- 0104
           ,x"4552" -- 0106
           ,x"5200" -- 0108
           ,x"0d0a" -- 010A
           ,x"434b" -- 010C
           ,x"534d" -- 010E
           ,x"2045" -- 0110
           ,x"5252" -- 0112
           ,x"000d" -- 0114
           ,x"0a54" -- 0116
           ,x"4147" -- 0118
           ,x"2045" -- 011A
           ,x"5252" -- 011C
           ,x"0055" -- 011E
           ,x"504c" -- 0120
           ,x"4420" -- 0122
           ,x"4552" -- 0124
           ,x"5200" -- 0126
           ,x"460d" -- 0128
           ,x"000a" -- 012A
           ,x"7f3a" -- 012C
           ,x"0d0a" -- 012E
           ,x"7f13" -- 0130
           ,x"0d14" -- 0132
           ,x"7f00" -- 0134
           ,x"120a" -- 0136
           ,x"7f00" -- 0138
           ,x"6242" -- 013A
           ,x"1100" -- 013C
           ,x"0000" -- 013E
           ,x"0400" -- 0140
           ,x"02e0" -- 0142
           ,x"ec00" -- 0144
           ,x"04c1" -- 0146
           ,x"0202" -- 0148
           ,x"fffc" -- 014A
           ,x"ccb1" -- 014C
           ,x"0201" -- 014E
           ,x"042e" -- 0150
           ,x"cc81" -- 0152
           ,x"0209" -- 0154
           ,x"0142" -- 0156
           ,x"04c1" -- 0158
           ,x"0641" -- 015A
           ,x"16fe" -- 015C
           ,x"c320" -- 015E
           ,x"013e" -- 0160
           ,x"c80c" -- 0162
           ,x"ec2e" -- 0164
           ,x"1f15" -- 0166
           ,x"1601" -- 0168
           ,x"2f45" -- 016A
           ,x"2fa0" -- 016C
           ,x"0014" -- 016E
           ,x"04c0" -- 0170
           ,x"0202" -- 0172
           ,x"0a05" -- 0174
           ,x"0203" -- 0176
           ,x"0004" -- 0178
           ,x"04c4" -- 017A
           ,x"0208" -- 017C
           ,x"0001" -- 017E
           ,x"2ec5" -- 0180
           ,x"0285" -- 0182
           ,x"0d00" -- 0184
           ,x"1604" -- 0186
           ,x"0205" -- 0188
           ,x"0a00" -- 018A
           ,x"2f05" -- 018C
           ,x"1019" -- 018E
           ,x"0285" -- 0190
           ,x"2000" -- 0192
           ,x"1316" -- 0194
           ,x"0285" -- 0196
           ,x"2c00" -- 0198
           ,x"1313" -- 019A
           ,x"0285" -- 019C
           ,x"4100" -- 019E
           ,x"113c" -- 01A0
           ,x"0285" -- 01A2
           ,x"5a00" -- 01A4
           ,x"1539" -- 01A6
           ,x"0603" -- 01A8
           ,x"1337" -- 01AA
           ,x"06c5" -- 01AC
           ,x"0245" -- 01AE
           ,x"001f" -- 01B0
           ,x"0283" -- 01B2
           ,x"0003" -- 01B4
           ,x"1301" -- 01B6
           ,x"0482" -- 01B8
           ,x"a105" -- 01BA
           ,x"0222" -- 01BC
           ,x"0050" -- 01BE
           ,x"10df" -- 01C0
           ,x"020b" -- 01C2
           ,x"027a" -- 01C4
           ,x"1002" -- 01C6
           ,x"022b" -- 01C8
           ,x"0004" -- 01CA
           ,x"c2bb" -- 01CC
           ,x"1325" -- 01CE
           ,x"810a" -- 01D0
           ,x"16fa" -- 01D2
           ,x"c1bb" -- 01D4
           ,x"c2db" -- 01D6
           ,x"0207" -- 01D8
           ,x"ec00" -- 01DA
           ,x"0285" -- 01DC
           ,x"0a00" -- 01DE
           ,x"130f" -- 01E0
           ,x"0916" -- 01E2
           ,x"170e" -- 01E4
           ,x"2e44" -- 01E6
           ,x"01f8" -- 01E8
           ,x"020e" -- 01EA
           ,x"cdc4" -- 01EC
           ,x"0583" -- 01EE
           ,x"0285" -- 01F0
           ,x"0d00" -- 01F2
           ,x"1306" -- 01F4
           ,x"10f5" -- 01F6
           ,x"05c7" -- 01F8
           ,x"0285" -- 01FA
           ,x"0d00" -- 01FC
           ,x"16f7" -- 01FE
           ,x"04c3" -- 0200
           ,x"045b" -- 0202
           ,x"04c0" -- 0204
           ,x"100b" -- 0206
           ,x"0200" -- 0208
           ,x"0001" -- 020A
           ,x"1008" -- 020C
           ,x"0200" -- 020E
           ,x"0002" -- 0210
           ,x"1005" -- 0212
           ,x"0200" -- 0214
           ,x"0003" -- 0216
           ,x"1002" -- 0218
           ,x"0200" -- 021A
           ,x"0004" -- 021C
           ,x"2fa0" -- 021E
           ,x"00a4" -- 0220
           ,x"2e00" -- 0222
           ,x"108e" -- 0224
           ,x"020c" -- 0226
           ,x"ec44" -- 0228
           ,x"04fc" -- 022A
           ,x"073c" -- 022C
           ,x"04fc" -- 022E
           ,x"04dc" -- 0230
           ,x"c320" -- 0232
           ,x"013e" -- 0234
           ,x"c80c" -- 0236
           ,x"ec2e" -- 0238
           ,x"1d1f" -- 023A
           ,x"04c3" -- 023C
           ,x"3220" -- 023E
           ,x"013a" -- 0240
           ,x"1e0d" -- 0242
           ,x"1f0f" -- 0244
           ,x"13fe" -- 0246
           ,x"0583" -- 0248
           ,x"1f0f" -- 024A
           ,x"16fd" -- 024C
           ,x"0207" -- 024E
           ,x"0084" -- 0250
           ,x"8dc3" -- 0252
           ,x"1102" -- 0254
           ,x"05c7" -- 0256
           ,x"10fc" -- 0258
           ,x"3317" -- 025A
           ,x"c1d7" -- 025C
           ,x"0287" -- 025E
           ,x"01a1" -- 0260
           ,x"1108" -- 0262
           ,x"1602" -- 0264
           ,x"0720" -- 0266
           ,x"ec44" -- 0268
           ,x"2f45" -- 026A
           ,x"0460" -- 026C
           ,x"1500" -- 026E
           ,x"0460" -- 0270
           ,x"0142" -- 0272
           ,x"05a0" -- 0274
           ,x"ec44" -- 0276
           ,x"10f8" -- 0278
           ,x"01a9" -- 027A
           ,x"0001" -- 027C
           ,x"036c" -- 027E
           ,x"01a4" -- 0280
           ,x"0003" -- 0282
           ,x"0334" -- 0284
           ,x"4ae9" -- 0286
           ,x"0001" -- 0288
           ,x"04ac" -- 028A
           ,x"0305" -- 028C
           ,x"0000" -- 028E
           ,x"042c" -- 0290
           ,x"0b05" -- 0292
           ,x"0001" -- 0294
           ,x"0436" -- 0296
           ,x"0273" -- 0298
           ,x"0000" -- 029A
           ,x"0426" -- 029C
           ,x"0dac" -- 029E
           ,x"0001" -- 02A0
           ,x"064a" -- 02A2
           ,x"0da4" -- 02A4
           ,x"0007" -- 02A6
           ,x"0552" -- 02A8
           ,x"0069" -- 02AA
           ,x"0003" -- 02AC
           ,x"0460" -- 02AE
           ,x"0249" -- 02B0
           ,x"0000" -- 02B2
           ,x"051a" -- 02B4
           ,x"0086" -- 02B6
           ,x"0007" -- 02B8
           ,x"0770" -- 02BA
           ,x"60a8" -- 02BC
           ,x"0003" -- 02BE
           ,x"07a0" -- 02C0
           ,x"19d4" -- 02C2
           ,x"0000" -- 02C4
           ,x"07b4" -- 02C6
           ,x"1438" -- 02C8
           ,x"0001" -- 02CA
           ,x"07c2" -- 02CC
           ,x"0038" -- 02CE
           ,x"0001" -- 02D0
           ,x"07ba" -- 02D2
           ,x"3078" -- 02D4
           ,x"0000" -- 02D6
           ,x"0e1a" -- 02D8
           ,x"0658" -- 02DA
           ,x"0003" -- 02DC
           ,x"1166" -- 02DE
           ,x"0000" -- 02E0
           ,x"1f15" -- 02E2
           ,x"16fe" -- 02E4
           ,x"04db" -- 02E6
           ,x"361b" -- 02E8
           ,x"1e12" -- 02EA
           ,x"0380" -- 02EC
           ,x"020a" -- 02EE
           ,x"186a" -- 02F0
           ,x"1d10" -- 02F2
           ,x"1f16" -- 02F4
           ,x"16fe" -- 02F6
           ,x"321b" -- 02F8
           ,x"d2db" -- 02FA
           ,x"0380" -- 02FC
           ,x"1000" -- 02FE
           ,x"160b" -- 0300
           ,x"c2e0" -- 0302
           ,x"ec44" -- 0304
           ,x"150e" -- 0306
           ,x"0a3a" -- 0308
           ,x"1f16" -- 030A
           ,x"16fe" -- 030C
           ,x"1f17" -- 030E
           ,x"16fc" -- 0310
           ,x"060a" -- 0312
           ,x"16fe" -- 0314
           ,x"0380" -- 0316
           ,x"c2e0" -- 0318
           ,x"ec46" -- 031A
           ,x"1303" -- 031C
           ,x"c2e0" -- 031E
           ,x"ec44" -- 0320
           ,x"11f3" -- 0322
           ,x"0380" -- 0324
           ,x"2f5b" -- 0326
           ,x"2f1b" -- 0328
           ,x"0380" -- 032A
           ,x"d33b" -- 032C
           ,x"13fd" -- 032E
           ,x"2f0c" -- 0330
           ,x"10fc" -- 0332
           ,x"4008" -- 0334
           ,x"4048" -- 0336
           ,x"0203" -- 0338
           ,x"0008" -- 033A
           ,x"2fa0" -- 033C
           ,x"00f2" -- 033E
           ,x"2e80" -- 0340
           ,x"2fa0" -- 0342
           ,x"00cf" -- 0344
           ,x"2e90" -- 0346
           ,x"1f15" -- 0348
           ,x"1602" -- 034A
           ,x"2f40" -- 034C
           ,x"0459" -- 034E
           ,x"8040" -- 0350
           ,x"13fd" -- 0352
           ,x"05c0" -- 0354
           ,x"0603" -- 0356
           ,x"0283" -- 0358
           ,x"0004" -- 035A
           ,x"1602" -- 035C
           ,x"2fa0" -- 035E
           ,x"0020" -- 0360
           ,x"c0c3" -- 0362
           ,x"13e9" -- 0364
           ,x"2fa0" -- 0366
           ,x"0020" -- 0368
           ,x"10ed" -- 036A
           ,x"4008" -- 036C
           ,x"1004" -- 036E
           ,x"0640" -- 0370
           ,x"0a25" -- 0372
           ,x"16fb" -- 0374
           ,x"8c30" -- 0376
           ,x"2fa0" -- 0378
           ,x"00f2" -- 037A
           ,x"2e80" -- 037C
           ,x"2fa0" -- 037E
           ,x"00cf" -- 0380
           ,x"2e90" -- 0382
           ,x"2fa0" -- 0384
           ,x"0020" -- 0386
           ,x"2e44" -- 0388
           ,x"0390" -- 038A
           ,x"020e" -- 038C
           ,x"c404" -- 038E
           ,x"0a25" -- 0390
           ,x"11ee" -- 0392
           ,x"0459" -- 0394
           ,x"04c9" -- 0396
           ,x"04cc" -- 0398
           ,x"2eca" -- 039A
           ,x"028a" -- 039C
           ,x"3000" -- 039E
           ,x"1a11" -- 03A0
           ,x"028a" -- 03A2
           ,x"3900" -- 03A4
           ,x"1208" -- 03A6
           ,x"028a" -- 03A8
           ,x"4100" -- 03AA
           ,x"1a0b" -- 03AC
           ,x"028a" -- 03AE
           ,x"4600" -- 03B0
           ,x"1b08" -- 03B2
           ,x"022a" -- 03B4
           ,x"0900" -- 03B6
           ,x"0a4a" -- 03B8
           ,x"09ca" -- 03BA
           ,x"0a4c" -- 03BC
           ,x"a30a" -- 03BE
           ,x"0589" -- 03C0
           ,x"10eb" -- 03C2
           ,x"028a" -- 03C4
           ,x"2000" -- 03C6
           ,x"130b" -- 03C8
           ,x"028a" -- 03CA
           ,x"2d00" -- 03CC
           ,x"1308" -- 03CE
           ,x"028a" -- 03D0
           ,x"0d00" -- 03D2
           ,x"1305" -- 03D4
           ,x"028a" -- 03D6
           ,x"2c00" -- 03D8
           ,x"160c" -- 03DA
           ,x"020a" -- 03DC
           ,x"2000" -- 03DE
           ,x"c249" -- 03E0
           ,x"1304" -- 03E2
           ,x"cecc" -- 03E4
           ,x"c6ca" -- 03E6
           ,x"8fbe" -- 03E8
           ,x"0380" -- 03EA
           ,x"05cb" -- 03EC
           ,x"c6ca" -- 03EE
           ,x"c39e" -- 03F0
           ,x"0380" -- 03F2
           ,x"05ce" -- 03F4
           ,x"10fc" -- 03F6
           ,x"c31b" -- 03F8
           ,x"0acc" -- 03FA
           ,x"0209" -- 03FC
           ,x"0001" -- 03FE
           ,x"1003" -- 0400
           ,x"c31b" -- 0402
           ,x"0209" -- 0404
           ,x"0004" -- 0406
           ,x"c28c" -- 0408
           ,x"09ca" -- 040A
           ,x"0a8a" -- 040C
           ,x"028a" -- 040E
           ,x"0900" -- 0410
           ,x"1202" -- 0412
           ,x"022a" -- 0414
           ,x"0700" -- 0416
           ,x"022a" -- 0418
           ,x"3000" -- 041A
           ,x"2f0a" -- 041C
           ,x"0bcc" -- 041E
           ,x"0609" -- 0420
           ,x"16f2" -- 0422
           ,x"0380" -- 0424
           ,x"0207" -- 0426
           ,x"9900" -- 0428
           ,x"03e0" -- 042A
           ,x"0380" -- 042C
           ,x"0287" -- 042E
           ,x"9900" -- 0430
           ,x"130b" -- 0432
           ,x"1013" -- 0434
           ,x"4008" -- 0436
           ,x"c190" -- 0438
           ,x"c420" -- 043A
           ,x"0440" -- 043C
           ,x"0380" -- 043E
           ,x"2fc0" -- 0440
           ,x"064e" -- 0442
           ,x"c406" -- 0444
           ,x"2fa0" -- 0446
           ,x"0023" -- 0448
           ,x"04c7" -- 044A
           ,x"020a" -- 044C
           ,x"fffa" -- 044E
           ,x"2fa0" -- 0450
           ,x"001e" -- 0452
           ,x"2eaa" -- 0454
           ,x"ec20" -- 0456
           ,x"05ca" -- 0458
           ,x"16fa" -- 045A
           ,x"0460" -- 045C
           ,x"0142" -- 045E
           ,x"c300" -- 0460
           ,x"04c7" -- 0462
           ,x"0241" -- 0464
           ,x"000f" -- 0466
           ,x"1303" -- 0468
           ,x"0281" -- 046A
           ,x"0009" -- 046C
           ,x"1a01" -- 046E
           ,x"0587" -- 0470
           ,x"0a61" -- 0472
           ,x"0208" -- 0474
           ,x"3406" -- 0476
           ,x"e201" -- 0478
           ,x"0488" -- 047A
           ,x"2fa0" -- 047C
           ,x"00f2" -- 047E
           ,x"2e8c" -- 0480
           ,x"2fa0" -- 0482
           ,x"00cf" -- 0484
           ,x"c1c7" -- 0486
           ,x"1601" -- 0488
           ,x"0986" -- 048A
           ,x"2e86" -- 048C
           ,x"2fa0" -- 048E
           ,x"0020" -- 0490
           ,x"2e44" -- 0492
           ,x"04a6" -- 0494
           ,x"020e" -- 0496
           ,x"c184" -- 0498
           ,x"c1c7" -- 049A
           ,x"1601" -- 049C
           ,x"0a86" -- 049E
           ,x"0248" -- 04A0
           ,x"f3ff" -- 04A2
           ,x"0488" -- 04A4
           ,x"09c5" -- 04A6
           ,x"16e5" -- 04A8
           ,x"0459" -- 04AA
           ,x"c1cd" -- 04AC
           ,x"c0c3" -- 04AE
           ,x"131f" -- 04B0
           ,x"0240" -- 04B2
           ,x"000f" -- 04B4
           ,x"c180" -- 04B6
           ,x"0a10" -- 04B8
           ,x"a1c0" -- 04BA
           ,x"2fa0" -- 04BC
           ,x"00bc" -- 04BE
           ,x"2e06" -- 04C0
           ,x"2fa0" -- 04C2
           ,x"00cf" -- 04C4
           ,x"2e97" -- 04C6
           ,x"2fa0" -- 04C8
           ,x"0020" -- 04CA
           ,x"2e44" -- 04CC
           ,x"04d4" -- 04CE
           ,x"020e" -- 04D0
           ,x"c5c4" -- 04D2
           ,x"0a25" -- 04D4
           ,x"153c" -- 04D6
           ,x"0a15" -- 04D8
           ,x"1304" -- 04DA
           ,x"0606" -- 04DC
           ,x"1138" -- 04DE
           ,x"0647" -- 04E0
           ,x"10ec" -- 04E2
           ,x"0286" -- 04E4
           ,x"000f" -- 04E6
           ,x"1333" -- 04E8
           ,x"0586" -- 04EA
           ,x"05c7" -- 04EC
           ,x"10e6" -- 04EE
           ,x"04c6" -- 04F0
           ,x"c1cd" -- 04F2
           ,x"2fa0" -- 04F4
           ,x"00bc" -- 04F6
           ,x"2e06" -- 04F8
           ,x"2fa0" -- 04FA
           ,x"00cf" -- 04FC
           ,x"2e97" -- 04FE
           ,x"0586" -- 0500
           ,x"05c7" -- 0502
           ,x"0286" -- 0504
           ,x"0008" -- 0506
           ,x"13f5" -- 0508
           ,x"0286" -- 050A
           ,x"0010" -- 050C
           ,x"1320" -- 050E
           ,x"2fa0" -- 0510
           ,x"0020" -- 0512
           ,x"2fa0" -- 0514
           ,x"00d6" -- 0516
           ,x"10ef" -- 0518
           ,x"0206" -- 051A
           ,x"003a" -- 051C
           ,x"0207" -- 051E
           ,x"0003" -- 0520
           ,x"0208" -- 0522
           ,x"ec1a" -- 0524
           ,x"2fa0" -- 0526
           ,x"00f2" -- 0528
           ,x"2f96" -- 052A
           ,x"2fa0" -- 052C
           ,x"00cf" -- 052E
           ,x"c118" -- 0530
           ,x"2e98" -- 0532
           ,x"2fa0" -- 0534
           ,x"0020" -- 0536
           ,x"2e44" -- 0538
           ,x"053e" -- 053A
           ,x"020e" -- 053C
           ,x"c604" -- 053E
           ,x"0a25" -- 0540
           ,x"1506" -- 0542
           ,x"0a15" -- 0544
           ,x"16ef" -- 0546
           ,x"05c6" -- 0548
           ,x"05c8" -- 054A
           ,x"0607" -- 054C
           ,x"16eb" -- 054E
           ,x"0459" -- 0550
           ,x"4008" -- 0552
           ,x"4048" -- 0554
           ,x"4088" -- 0556
           ,x"8040" -- 0558
           ,x"1202" -- 055A
           ,x"0460" -- 055C
           ,x"0214" -- 055E
           ,x"04c4" -- 0560
           ,x"04c3" -- 0562
           ,x"2fa0" -- 0564
           ,x"0028" -- 0566
           ,x"2f44" -- 0568
           ,x"0284" -- 056A
           ,x"0d00" -- 056C
           ,x"1603" -- 056E
           ,x"0204" -- 0570
           ,x"2000" -- 0572
           ,x"1001" -- 0574
           ,x"2f04" -- 0576
           ,x"d8c4" -- 0578
           ,x"ec0c" -- 057A
           ,x"0583" -- 057C
           ,x"0283" -- 057E
           ,x"0008" -- 0580
           ,x"1304" -- 0582
           ,x"0284" -- 0584
           ,x"2000" -- 0586
           ,x"16ef" -- 0588
           ,x"10f6" -- 058A
           ,x"2fa0" -- 058C
           ,x"002d" -- 058E
           ,x"2f44" -- 0590
           ,x"0284" -- 0592
           ,x"5900" -- 0594
           ,x"1641" -- 0596
           ,x"04e0" -- 0598
           ,x"ec46" -- 059A
           ,x"2fa0" -- 059C
           ,x"0136" -- 059E
           ,x"04ca" -- 05A0
           ,x"04c5" -- 05A2
           ,x"06a0" -- 05A4
           ,x"061c" -- 05A6
           ,x"3000" -- 05A8
           ,x"2fa0" -- 05AA
           ,x"ec0c" -- 05AC
           ,x"0203" -- 05AE
           ,x"0008" -- 05B0
           ,x"d123" -- 05B2
           ,x"ec0b" -- 05B4
           ,x"0984" -- 05B6
           ,x"a144" -- 05B8
           ,x"0603" -- 05BA
           ,x"16fa" -- 05BC
           ,x"c282" -- 05BE
           ,x"06a0" -- 05C0
           ,x"061c" -- 05C2
           ,x"3100" -- 05C4
           ,x"c280" -- 05C6
           ,x"06a0" -- 05C8
           ,x"061c" -- 05CA
           ,x"3900" -- 05CC
           ,x"c290" -- 05CE
           ,x"06a0" -- 05D0
           ,x"061c" -- 05D2
           ,x"4200" -- 05D4
           ,x"8040" -- 05D6
           ,x"1304" -- 05D8
           ,x"05c0" -- 05DA
           ,x"0283" -- 05DC
           ,x"003c" -- 05DE
           ,x"1af6" -- 05E0
           ,x"0225" -- 05E2
           ,x"0037" -- 05E4
           ,x"c285" -- 05E6
           ,x"050a" -- 05E8
           ,x"06a0" -- 05EA
           ,x"061c" -- 05EC
           ,x"3700" -- 05EE
           ,x"04c5" -- 05F0
           ,x"2fa0" -- 05F2
           ,x"0128" -- 05F4
           ,x"8040" -- 05F6
           ,x"1304" -- 05F8
           ,x"04c3" -- 05FA
           ,x"2fa0" -- 05FC
           ,x"0137" -- 05FE
           ,x"10e2" -- 0600
           ,x"2fa0" -- 0602
           ,x"012b" -- 0604
           ,x"0203" -- 0606
           ,x"003c" -- 0608
           ,x"2fa0" -- 060A
           ,x"0134" -- 060C
           ,x"0603" -- 060E
           ,x"16fc" -- 0610
           ,x"0720" -- 0612
           ,x"ec46" -- 0614
           ,x"2fa0" -- 0616
           ,x"00f2" -- 0618
           ,x"104a" -- 061A
           ,x"c13b" -- 061C
           ,x"2f04" -- 061E
           ,x"0984" -- 0620
           ,x"a144" -- 0622
           ,x"2e8a" -- 0624
           ,x"0223" -- 0626
           ,x"0005" -- 0628
           ,x"0204" -- 062A
           ,x"0004" -- 062C
           ,x"0b4a" -- 062E
           ,x"c30a" -- 0630
           ,x"09cc" -- 0632
           ,x"a14c" -- 0634
           ,x"0225" -- 0636
           ,x"0030" -- 0638
           ,x"028c" -- 063A
           ,x"000a" -- 063C
           ,x"1a02" -- 063E
           ,x"0225" -- 0640
           ,x"0007" -- 0642
           ,x"0604" -- 0644
           ,x"16f3" -- 0646
           ,x"045b" -- 0648
           ,x"2fa0" -- 064A
           ,x"002d" -- 064C
           ,x"2f44" -- 064E
           ,x"0284" -- 0650
           ,x"5900" -- 0652
           ,x"162d" -- 0654
           ,x"0206" -- 0656
           ,x"1100" -- 0658
           ,x"2f06" -- 065A
           ,x"04c7" -- 065C
           ,x"04c8" -- 065E
           ,x"06a0" -- 0660
           ,x"0728" -- 0662
           ,x"100b" -- 0664
           ,x"d22a" -- 0666
           ,x"070e" -- 0668
           ,x"132d" -- 066A
           ,x"06a0" -- 066C
           ,x"0722" -- 066E
           ,x"100e" -- 0670
           ,x"0205" -- 0672
           ,x"0008" -- 0674
           ,x"0878" -- 0676
           ,x"0468" -- 0678
           ,x"0678" -- 067A
           ,x"0286" -- 067C
           ,x"0047" -- 067E
           ,x"1106" -- 0680
           ,x"0286" -- 0682
           ,x"004a" -- 0684
           ,x"1516" -- 0686
           ,x"0226" -- 0688
           ,x"ffc9" -- 068A
           ,x"10ec" -- 068C
           ,x"0286" -- 068E
           ,x"003a" -- 0690
           ,x"1610" -- 0692
           ,x"04ca" -- 0694
           ,x"0705" -- 0696
           ,x"020c" -- 0698
           ,x"0080" -- 069A
           ,x"1f0f" -- 069C
           ,x"16fb" -- 069E
           ,x"0605" -- 06A0
           ,x"16fc" -- 06A2
           ,x"c28a" -- 06A4
           ,x"1609" -- 06A6
           ,x"2fa0" -- 06A8
           ,x"00f2" -- 06AA
           ,x"2fa0" -- 06AC
           ,x"ec02" -- 06AE
           ,x"0460" -- 06B0
           ,x"0142" -- 06B2
           ,x"04c0" -- 06B4
           ,x"070a" -- 06B6
           ,x"10ee" -- 06B8
           ,x"c000" -- 06BA
           ,x"1302" -- 06BC
           ,x"0460" -- 06BE
           ,x"0208" -- 06C0
           ,x"0460" -- 06C2
           ,x"0204" -- 06C4
           ,x"2f46" -- 06C6
           ,x"9806" -- 06C8
           ,x"00f2" -- 06CA
           ,x"16fc" -- 06CC
           ,x"10c6" -- 06CE
           ,x"a280" -- 06D0
           ,x"c24a" -- 06D2
           ,x"10c4" -- 06D4
           ,x"a280" -- 06D6
           ,x"ce4a" -- 06D8
           ,x"10c1" -- 06DA
           ,x"a1ca" -- 06DC
           ,x"13bf" -- 06DE
           ,x"0200" -- 06E0
           ,x"0001" -- 06E2
           ,x"10e8" -- 06E4
           ,x"020a" -- 06E6
           ,x"ec02" -- 06E8
           ,x"1003" -- 06EA
           ,x"0645" -- 06EC
           ,x"020a" -- 06EE
           ,x"ec22" -- 06F0
           ,x"2f46" -- 06F2
           ,x"de86" -- 06F4
           ,x"0986" -- 06F6
           ,x"a1c6" -- 06F8
           ,x"0605" -- 06FA
           ,x"16fa" -- 06FC
           ,x"10af" -- 06FE
           ,x"a280" -- 0700
           ,x"c38a" -- 0702
           ,x"10ac" -- 0704
           ,x"024a" -- 0706
           ,x"fffe" -- 0708
           ,x"c00a" -- 070A
           ,x"10a8" -- 070C
           ,x"3745" -- 070E
           ,x"443a" -- 0710
           ,x"3a3a" -- 0712
           ,x"3a32" -- 0714
           ,x"f22d" -- 0716
           ,x"2c30" -- 0718
           ,x"2f47" -- 071A
           ,x"1e00" -- 071C
           ,x"3a3a" -- 071E
           ,x"3bf3" -- 0720
           ,x"0205" -- 0722
           ,x"fffc" -- 0724
           ,x"1001" -- 0726
           ,x"0705" -- 0728
           ,x"04ca" -- 072A
           ,x"2f46" -- 072C
           ,x"0286" -- 072E
           ,x"2000" -- 0730
           ,x"11fc" -- 0732
           ,x"0286" -- 0734
           ,x"5f00" -- 0736
           ,x"15f9" -- 0738
           ,x"0986" -- 073A
           ,x"0288" -- 073C
           ,x"3200" -- 073E
           ,x"1301" -- 0740
           ,x"a1c6" -- 0742
           ,x"0286" -- 0744
           ,x"0030" -- 0746
           ,x"1112" -- 0748
           ,x"0286" -- 074A
           ,x"0039" -- 074C
           ,x"1208" -- 074E
           ,x"0286" -- 0750
           ,x"0041" -- 0752
           ,x"110c" -- 0754
           ,x"0286" -- 0756
           ,x"0046" -- 0758
           ,x"1509" -- 075A
           ,x"0226" -- 075C
           ,x"0009" -- 075E
           ,x"0246" -- 0760
           ,x"000f" -- 0762
           ,x"0a4a" -- 0764
           ,x"a286" -- 0766
           ,x"0585" -- 0768
           ,x"16e0" -- 076A
           ,x"05cb" -- 076C
           ,x"045b" -- 076E
           ,x"0203" -- 0770
           ,x"8402" -- 0772
           ,x"0204" -- 0774
           ,x"05c0" -- 0776
           ,x"0a25" -- 0778
           ,x"1103" -- 077A
           ,x"4008" -- 077C
           ,x"4048" -- 077E
           ,x"1007" -- 0780
           ,x"0223" -- 0782
           ,x"1000" -- 0784
           ,x"0224" -- 0786
           ,x"ffc0" -- 0788
           ,x"0a82" -- 078A
           ,x"1001" -- 078C
           ,x"0484" -- 078E
           ,x"0483" -- 0790
           ,x"1603" -- 0792
           ,x"2fa0" -- 0794
           ,x"00f2" -- 0796
           ,x"2e80" -- 0798
           ,x"8040" -- 079A
           ,x"16f8" -- 079C
           ,x"0459" -- 079E
           ,x"2fa0" -- 07A0
           ,x"00c0" -- 07A2
           ,x"c100" -- 07A4
           ,x"a101" -- 07A6
           ,x"2e84" -- 07A8
           ,x"2fa0" -- 07AA
           ,x"00c9" -- 07AC
           ,x"6001" -- 07AE
           ,x"2e80" -- 07B0
           ,x"0459" -- 07B2
           ,x"0560" -- 07B4
           ,x"ec44" -- 07B6
           ,x"0459" -- 07B8
           ,x"04e0" -- 07BA
           ,x"ec4e" -- 07BC
           ,x"04e0" -- 07BE
           ,x"ec4c" -- 07C0
           ,x"c240" -- 07C2
           ,x"2fa0" -- 07C4
           ,x"00f2" -- 07C6
           ,x"020a" -- 07C8
           ,x"0850" -- 07CA
           ,x"0200" -- 07CC
           ,x"ec52" -- 07CE
           ,x"0208" -- 07D0
           ,x"0006" -- 07D2
           ,x"04f0" -- 07D4
           ,x"0608" -- 07D6
           ,x"15fd" -- 07D8
           ,x"2e89" -- 07DA
           ,x"2fa0" -- 07DC
           ,x"001c" -- 07DE
           ,x"069a" -- 07E0
           ,x"0284" -- 07E2
           ,x"0020" -- 07E4
           ,x"1316" -- 07E6
           ,x"0284" -- 07E8
           ,x"002a" -- 07EA
           ,x"1605" -- 07EC
           ,x"069a" -- 07EE
           ,x"0284" -- 07F0
           ,x"000d" -- 07F2
           ,x"16fc" -- 07F4
           ,x"10e6" -- 07F6
           ,x"06a0" -- 07F8
           ,x"0bee" -- 07FA
           ,x"c807" -- 07FC
           ,x"ec52" -- 07FE
           ,x"c809" -- 0800
           ,x"ec54" -- 0802
           ,x"c107" -- 0804
           ,x"06a0" -- 0806
           ,x"0c64" -- 0808
           ,x"1321" -- 080A
           ,x"9807" -- 080C
           ,x"0bf3" -- 080E
           ,x"1303" -- 0810
           ,x"1004" -- 0812
           ,x"2fa0" -- 0814
           ,x"0021" -- 0816
           ,x"2fa0" -- 0818
           ,x"0021" -- 081A
           ,x"0207" -- 081C
           ,x"0ce3" -- 081E
           ,x"04c5" -- 0820
           ,x"04c6" -- 0822
           ,x"069a" -- 0824
           ,x"06a0" -- 0826
           ,x"0c34" -- 0828
           ,x"1643" -- 082A
           ,x"0ab4" -- 082C
           ,x"0587" -- 082E
           ,x"d017" -- 0830
           ,x"1102" -- 0832
           ,x"1372" -- 0834
           ,x"05c6" -- 0836
           ,x"0a10" -- 0838
           ,x"09e0" -- 083A
           ,x"8005" -- 083C
           ,x"11f7" -- 083E
           ,x"156c" -- 0840
           ,x"d017" -- 0842
           ,x"0a30" -- 0844
           ,x"9100" -- 0846
           ,x"16f2" -- 0848
           ,x"0585" -- 084A
           ,x"10eb" -- 084C
           ,x"1065" -- 084E
           ,x"2f44" -- 0850
           ,x"0284" -- 0852
           ,x"1b00" -- 0854
           ,x"13b6" -- 0856
           ,x"0284" -- 0858
           ,x"2000" -- 085A
           ,x"1a01" -- 085C
           ,x"2f04" -- 085E
           ,x"0984" -- 0860
           ,x"c804" -- 0862
           ,x"ec60" -- 0864
           ,x"045b" -- 0866
           ,x"069a" -- 0868
           ,x"0284" -- 086A
           ,x"0027" -- 086C
           ,x"1655" -- 086E
           ,x"c1c9" -- 0870
           ,x"75d7" -- 0872
           ,x"0588" -- 0874
           ,x"069a" -- 0876
           ,x"0284" -- 0878
           ,x"0027" -- 087A
           ,x"1358" -- 087C
           ,x"06c4" -- 087E
           ,x"ddc4" -- 0880
           ,x"10f7" -- 0882
           ,x"06a0" -- 0884
           ,x"0b14" -- 0886
           ,x"c806" -- 0888
           ,x"ec54" -- 088A
           ,x"1064" -- 088C
           ,x"070e" -- 088E
           ,x"c006" -- 0890
           ,x"06a0" -- 0892
           ,x"0b14" -- 0894
           ,x"c809" -- 0896
           ,x"ec54" -- 0898
           ,x"0280" -- 089A
           ,x"0014" -- 089C
           ,x"1605" -- 089E
           ,x"a189" -- 08A0
           ,x"1303" -- 08A2
           ,x"0586" -- 08A4
           ,x"8246" -- 08A6
           ,x"1a38" -- 08A8
           ,x"c246" -- 08AA
           ,x"0249" -- 08AC
           ,x"fffe" -- 08AE
           ,x"1052" -- 08B0
           ,x"c145" -- 08B2
           ,x"13af" -- 08B4
           ,x"d017" -- 08B6
           ,x"1130" -- 08B8
           ,x"070e" -- 08BA
           ,x"0286" -- 08BC
           ,x"0032" -- 08BE
           ,x"13e1" -- 08C0
           ,x"0286" -- 08C2
           ,x"009a" -- 08C4
           ,x"13d0" -- 08C6
           ,x"c026" -- 08C8
           ,x"0d76" -- 08CA
           ,x"c040" -- 08CC
           ,x"0241" -- 08CE
           ,x"fff0" -- 08D0
           ,x"1302" -- 08D2
           ,x"c641" -- 08D4
           ,x"05c8" -- 08D6
           ,x"c040" -- 08D8
           ,x"0241" -- 08DA
           ,x"000f" -- 08DC
           ,x"d021" -- 08DE
           ,x"0cd6" -- 08E0
           ,x"06c0" -- 08E2
           ,x"0260" -- 08E4
           ,x"ffe0" -- 08E6
           ,x"c040" -- 08E8
           ,x"0921" -- 08EA
           ,x"0241" -- 08EC
           ,x"0006" -- 08EE
           ,x"c061" -- 08F0
           ,x"0cc6" -- 08F2
           ,x"1307" -- 08F4
           ,x"0284" -- 08F6
           ,x"0020" -- 08F8
           ,x"160f" -- 08FA
           ,x"04ce" -- 08FC
           ,x"020f" -- 08FE
           ,x"0904" -- 0900
           ,x"0691" -- 0902
           ,x"c040" -- 0904
           ,x"0ad1" -- 0906
           ,x"09c1" -- 0908
           ,x"c061" -- 090A
           ,x"0cc6" -- 090C
           ,x"1309" -- 090E
           ,x"04c0" -- 0910
           ,x"04ce" -- 0912
           ,x"020f" -- 0914
           ,x"0922" -- 0916
           ,x"0691" -- 0918
           ,x"2fa0" -- 091A
           ,x"00d1" -- 091C
           ,x"0460" -- 091E
           ,x"07c4" -- 0920
           ,x"0284" -- 0922
           ,x"000d" -- 0924
           ,x"1307" -- 0926
           ,x"0284" -- 0928
           ,x"0020" -- 092A
           ,x"16f6" -- 092C
           ,x"069a" -- 092E
           ,x"0284" -- 0930
           ,x"000d" -- 0932
           ,x"16fc" -- 0934
           ,x"0280" -- 0936
           ,x"0030" -- 0938
           ,x"135c" -- 093A
           ,x"2f20" -- 093C
           ,x"00f2" -- 093E
           ,x"2e89" -- 0940
           ,x"c089" -- 0942
           ,x"06a0" -- 0944
           ,x"0c86" -- 0946
           ,x"0204" -- 0948
           ,x"2052" -- 094A
           ,x"c0c3" -- 094C
           ,x"1301" -- 094E
           ,x"06c4" -- 0950
           ,x"2f04" -- 0952
           ,x"2eb9" -- 0954
           ,x"2fa0" -- 0956
           ,x"00f2" -- 0958
           ,x"0648" -- 095A
           ,x"15f1" -- 095C
           ,x"0200" -- 095E
           ,x"ec56" -- 0960
           ,x"06a0" -- 0962
           ,x"0c9a" -- 0964
           ,x"06a0" -- 0966
           ,x"0c9a" -- 0968
           ,x"c120" -- 096A
           ,x"ec52" -- 096C
           ,x"1331" -- 096E
           ,x"0224" -- 0970
           ,x"8000" -- 0972
           ,x"06a0" -- 0974
           ,x"0c64" -- 0976
           ,x"1608" -- 0978
           ,x"06a0" -- 097A
           ,x"09d6" -- 097C
           ,x"c390" -- 097E
           ,x"c403" -- 0980
           ,x"06a0" -- 0982
           ,x"09e6" -- 0984
           ,x"c00e" -- 0986
           ,x"16fa" -- 0988
           ,x"0224" -- 098A
           ,x"8080" -- 098C
           ,x"06a0" -- 098E
           ,x"0c64" -- 0990
           ,x"161a" -- 0992
           ,x"06a0" -- 0994
           ,x"09d6" -- 0996
           ,x"04ce" -- 0998
           ,x"0580" -- 099A
           ,x"d390" -- 099C
           ,x"c083" -- 099E
           ,x"6080" -- 09A0
           ,x"0602" -- 09A2
           ,x"0a72" -- 09A4
           ,x"1907" -- 09A6
           ,x"0600" -- 09A8
           ,x"2e80" -- 09AA
           ,x"2fa0" -- 09AC
           ,x"00d1" -- 09AE
           ,x"2fa0" -- 09B0
           ,x"00f2" -- 09B2
           ,x"1004" -- 09B4
           ,x"d402" -- 09B6
           ,x"0600" -- 09B8
           ,x"06a0" -- 09BA
           ,x"09e6" -- 09BC
           ,x"087e" -- 09BE
           ,x"05ce" -- 09C0
           ,x"1302" -- 09C2
           ,x"a00e" -- 09C4
           ,x"10e8" -- 09C6
           ,x"0200" -- 09C8
           ,x"ec52" -- 09CA
           ,x"04c4" -- 09CC
           ,x"06a0" -- 09CE
           ,x"0c9c" -- 09D0
           ,x"0460" -- 09D2
           ,x"07c8" -- 09D4
           ,x"c012" -- 09D6
           ,x"04e2" -- 09D8
           ,x"fffe" -- 09DA
           ,x"0620" -- 09DC
           ,x"ec4c" -- 09DE
           ,x"c0e0" -- 09E0
           ,x"ec54" -- 09E2
           ,x"045b" -- 09E4
           ,x"2e80" -- 09E6
           ,x"2f20" -- 09E8
           ,x"0a05" -- 09EA
           ,x"2e90" -- 09EC
           ,x"2fa0" -- 09EE
           ,x"00f2" -- 09F0
           ,x"045b" -- 09F2
           ,x"2fa0" -- 09F4
           ,x"001f" -- 09F6
           ,x"2ea0" -- 09F8
           ,x"ec4c" -- 09FA
           ,x"0460" -- 09FC
           ,x"0142" -- 09FE
           ,x"069a" -- 0A00
           ,x"0284" -- 0A02
           ,x"002a" -- 0A04
           ,x"131a" -- 0A06
           ,x"0284" -- 0A08
           ,x"0040" -- 0A0A
           ,x"1622" -- 0A0C
           ,x"06a0" -- 0A0E
           ,x"0b14" -- 0A10
           ,x"c088" -- 0A12
           ,x"a089" -- 0A14
           ,x"c486" -- 0A16
           ,x"05c8" -- 0A18
           ,x"0206" -- 0A1A
           ,x"0020" -- 0A1C
           ,x"0284" -- 0A1E
           ,x"0028" -- 0A20
           ,x"1608" -- 0A22
           ,x"06a0" -- 0A24
           ,x"0ad0" -- 0A26
           ,x"0266" -- 0A28
           ,x"0020" -- 0A2A
           ,x"0284" -- 0A2C
           ,x"0029" -- 0A2E
           ,x"1649" -- 0A30
           ,x"069a" -- 0A32
           ,x"c000" -- 0A34
           ,x"1601" -- 0A36
           ,x"0a66" -- 0A38
           ,x"1040" -- 0A3A
           ,x"06a0" -- 0A3C
           ,x"0ad0" -- 0A3E
           ,x"0266" -- 0A40
           ,x"0010" -- 0A42
           ,x"0284" -- 0A44
           ,x"002b" -- 0A46
           ,x"1603" -- 0A48
           ,x"069a" -- 0A4A
           ,x"0266" -- 0A4C
           ,x"0030" -- 0A4E
           ,x"10f1" -- 0A50
           ,x"020e" -- 0A52
           ,x"0a34" -- 0A54
           ,x"c80e" -- 0A56
           ,x"ec5e" -- 0A58
           ,x"0460" -- 0A5A
           ,x"0ad6" -- 0A5C
           ,x"06a0" -- 0A5E
           ,x"0ad0" -- 0A60
           ,x"0a46" -- 0A62
           ,x"102b" -- 0A64
           ,x"c006" -- 0A66
           ,x"0280" -- 0A68
           ,x"0030" -- 0A6A
           ,x"1604" -- 0A6C
           ,x"0284" -- 0A6E
           ,x"000d" -- 0A70
           ,x"1312" -- 0A72
           ,x"070e" -- 0A74
           ,x"06a0" -- 0A76
           ,x"0b14" -- 0A78
           ,x"0280" -- 0A7A
           ,x"0030" -- 0A7C
           ,x"130b" -- 0A7E
           ,x"c089" -- 0A80
           ,x"a088" -- 0A82
           ,x"c486" -- 0A84
           ,x"05c8" -- 0A86
           ,x"0280" -- 0A88
           ,x"0026" -- 0A8A
           ,x"1605" -- 0A8C
           ,x"070e" -- 0A8E
           ,x"0284" -- 0A90
           ,x"002c" -- 0A92
           ,x"13f0" -- 0A94
           ,x"c386" -- 0A96
           ,x"045f" -- 0A98
           ,x"06a0" -- 0A9A
           ,x"0ad0" -- 0A9C
           ,x"10ca" -- 0A9E
           ,x"06a0" -- 0AA0
           ,x"0b14" -- 0AA2
           ,x"c089" -- 0AA4
           ,x"05c2" -- 0AA6
           ,x"6182" -- 0AA8
           ,x"0816" -- 0AAA
           ,x"0286" -- 0AAC
           ,x"007f" -- 0AAE
           ,x"1507" -- 0AB0
           ,x"0286" -- 0AB2
           ,x"ff80" -- 0AB4
           ,x"1104" -- 0AB6
           ,x"0246" -- 0AB8
           ,x"00ff" -- 0ABA
           ,x"e646" -- 0ABC
           ,x"045f" -- 0ABE
           ,x"2fa0" -- 0AC0
           ,x"00d6" -- 0AC2
           ,x"0460" -- 0AC4
           ,x"091a" -- 0AC6
           ,x"070e" -- 0AC8
           ,x"06a0" -- 0ACA
           ,x"0b14" -- 0ACC
           ,x"10ee" -- 0ACE
           ,x"c80b" -- 0AD0
           ,x"ec5e" -- 0AD2
           ,x"069a" -- 0AD4
           ,x"020c" -- 0AD6
           ,x"0b04" -- 0AD8
           ,x"0284" -- 0ADA
           ,x"0052" -- 0ADC
           ,x"130c" -- 0ADE
           ,x"0284" -- 0AE0
           ,x"003a" -- 0AE2
           ,x"110a" -- 0AE4
           ,x"0284" -- 0AE6
           ,x"003e" -- 0AE8
           ,x"1309" -- 0AEA
           ,x"020e" -- 0AEC
           ,x"fffe" -- 0AEE
           ,x"020d" -- 0AF0
           ,x"0b04" -- 0AF2
           ,x"0460" -- 0AF4
           ,x"0b18" -- 0AF6
           ,x"069a" -- 0AF8
           ,x"0460" -- 0AFA
           ,x"0c2a" -- 0AFC
           ,x"069a" -- 0AFE
           ,x"0460" -- 0B00
           ,x"0c0c" -- 0B02
           ,x"c145" -- 0B04
           ,x"11de" -- 0B06
           ,x"0286" -- 0B08
           ,x"0010" -- 0B0A
           ,x"14db" -- 0B0C
           ,x"c2e0" -- 0B0E
           ,x"ec5e" -- 0B10
           ,x"045b" -- 0B12
           ,x"c34b" -- 0B14
           ,x"069a" -- 0B16
           ,x"04e0" -- 0B18
           ,x"ec50" -- 0B1A
           ,x"0284" -- 0B1C
           ,x"0027" -- 0B1E
           ,x"1307" -- 0B20
           ,x"0284" -- 0B22
           ,x"002d" -- 0B24
           ,x"1610" -- 0B26
           ,x"054d" -- 0B28
           ,x"05ce" -- 0B2A
           ,x"069a" -- 0B2C
           ,x"1011" -- 0B2E
           ,x"04c6" -- 0B30
           ,x"04ce" -- 0B32
           ,x"069a" -- 0B34
           ,x"0284" -- 0B36
           ,x"0027" -- 0B38
           ,x"1304" -- 0B3A
           ,x"06c6" -- 0B3C
           ,x"d106" -- 0B3E
           ,x"c184" -- 0B40
           ,x"10f8" -- 0B42
           ,x"069a" -- 0B44
           ,x"1043" -- 0B46
           ,x"0284" -- 0B48
           ,x"002b" -- 0B4A
           ,x"13ee" -- 0B4C
           ,x"c38e" -- 0B4E
           ,x"154b" -- 0B50
           ,x"0284" -- 0B52
           ,x"0024" -- 0B54
           ,x"1603" -- 0B56
           ,x"c189" -- 0B58
           ,x"069a" -- 0B5A
           ,x"1037" -- 0B5C
           ,x"0284" -- 0B5E
           ,x"003e" -- 0B60
           ,x"1604" -- 0B62
           ,x"069a" -- 0B64
           ,x"06a0" -- 0B66
           ,x"0c0a" -- 0B68
           ,x"1030" -- 0B6A
           ,x"06a0" -- 0B6C
           ,x"0c34" -- 0B6E
           ,x"11a9" -- 0B70
           ,x"1325" -- 0B72
           ,x"06a0" -- 0B74
           ,x"0c28" -- 0B76
           ,x"1029" -- 0B78
           ,x"c38e" -- 0B7A
           ,x"16a3" -- 0B7C
           ,x"c059" -- 0B7E
           ,x"04c2" -- 0B80
           ,x"06a0" -- 0B82
           ,x"0c86" -- 0B84
           ,x"c4c9" -- 0B86
           ,x"0241" -- 0B88
           ,x"f000" -- 0B8A
           ,x"0281" -- 0B8C
           ,x"1000" -- 0B8E
           ,x"1611" -- 0B90
           ,x"0264" -- 0B92
           ,x"0080" -- 0B94
           ,x"c189" -- 0B96
           ,x"0643" -- 0B98
           ,x"c4c4" -- 0B9A
           ,x"8820" -- 0B9C
           ,x"ec56" -- 0B9E
           ,x"ec5a" -- 0BA0
           ,x"1603" -- 0BA2
           ,x"c1a0" -- 0BA4
           ,x"ec58" -- 0BA6
           ,x"1012" -- 0BA8
           ,x"06a0" -- 0BAA
           ,x"0c64" -- 0BAC
           ,x"1601" -- 0BAE
           ,x"c192" -- 0BB0
           ,x"100d" -- 0BB2
           ,x"a4c8" -- 0BB4
           ,x"0264" -- 0BB6
           ,x"8000" -- 0BB8
           ,x"04c6" -- 0BBA
           ,x"10ed" -- 0BBC
           ,x"06a0" -- 0BBE
           ,x"0bee" -- 0BC0
           ,x"c107" -- 0BC2
           ,x"06a0" -- 0BC4
           ,x"0c64" -- 0BC6
           ,x"16d8" -- 0BC8
           ,x"c192" -- 0BCA
           ,x"05ce" -- 0BCC
           ,x"c120" -- 0BCE
           ,x"ec60" -- 0BD0
           ,x"c34d" -- 0BD2
           ,x"1502" -- 0BD4
           ,x"0506" -- 0BD6
           ,x"054d" -- 0BD8
           ,x"c145" -- 0BDA
           ,x"1194" -- 0BDC
           ,x"c38e" -- 0BDE
           ,x"1305" -- 0BE0
           ,x"a806" -- 0BE2
           ,x"ec50" -- 0BE4
           ,x"109d" -- 0BE6
           ,x"c1a0" -- 0BE8
           ,x"ec50" -- 0BEA
           ,x"045d" -- 0BEC
           ,x"c30b" -- 0BEE
           ,x"0207" -- 0BF0
           ,x"0031" -- 0BF2
           ,x"06a0" -- 0BF4
           ,x"0c34" -- 0BF6
           ,x"111c" -- 0BF8
           ,x"1303" -- 0BFA
           ,x"0a87" -- 0BFC
           ,x"1919" -- 0BFE
           ,x"1001" -- 0C00
           ,x"0a87" -- 0C02
           ,x"a1c4" -- 0C04
           ,x"069a" -- 0C06
           ,x"10f5" -- 0C08
           ,x"c30b" -- 0C0A
           ,x"0202" -- 0C0C
           ,x"0010" -- 0C0E
           ,x"04c6" -- 0C10
           ,x"0705" -- 0C12
           ,x"06a0" -- 0C14
           ,x"0c34" -- 0C16
           ,x"110c" -- 0C18
           ,x"8083" -- 0C1A
           ,x"1409" -- 0C1C
           ,x"c146" -- 0C1E
           ,x"3942" -- 0C20
           ,x"a183" -- 0C22
           ,x"069a" -- 0C24
           ,x"10f6" -- 0C26
           ,x"c30b" -- 0C28
           ,x"0202" -- 0C2A
           ,x"000a" -- 0C2C
           ,x"10f0" -- 0C2E
           ,x"0705" -- 0C30
           ,x"045c" -- 0C32
           ,x"0701" -- 0C34
           ,x"c0c4" -- 0C36
           ,x"0284" -- 0C38
           ,x"0024" -- 0C3A
           ,x"1306" -- 0C3C
           ,x"0223" -- 0C3E
           ,x"ffd0" -- 0C40
           ,x"170e" -- 0C42
           ,x"0283" -- 0C44
           ,x"0009" -- 0C46
           ,x"1502" -- 0C48
           ,x"0501" -- 0C4A
           ,x"045b" -- 0C4C
           ,x"0223" -- 0C4E
           ,x"fff9" -- 0C50
           ,x"0283" -- 0C52
           ,x"000a" -- 0C54
           ,x"1a04" -- 0C56
           ,x"0283" -- 0C58
           ,x"0023" -- 0C5A
           ,x"1b01" -- 0C5C
           ,x"04c1" -- 0C5E
           ,x"c041" -- 0C60
           ,x"045b" -- 0C62
           ,x"0703" -- 0C64
           ,x"c060" -- 0C66
           ,x"ec4e" -- 0C68
           ,x"130b" -- 0C6A
           ,x"0a21" -- 0C6C
           ,x"0202" -- 0C6E
           ,x"ec62" -- 0C70
           ,x"a042" -- 0C72
           ,x"04c3" -- 0C74
           ,x"05c2" -- 0C76
           ,x"8c84" -- 0C78
           ,x"1303" -- 0C7A
           ,x"8042" -- 0C7C
           ,x"1afb" -- 0C7E
           ,x"0583" -- 0C80
           ,x"c0c3" -- 0C82
           ,x"045b" -- 0C84
           ,x"0203" -- 0C86
           ,x"ec58" -- 0C88
           ,x"84c2" -- 0C8A
           ,x"1305" -- 0C8C
           ,x"0203" -- 0C8E
           ,x"ec5c" -- 0C90
           ,x"84c2" -- 0C92
           ,x"1301" -- 0C94
           ,x"04c3" -- 0C96
           ,x"045b" -- 0C98
           ,x"c110" -- 0C9A
           ,x"c30b" -- 0C9C
           ,x"06a0" -- 0C9E
           ,x"0c64" -- 0CA0
           ,x"130d" -- 0CA2
           ,x"c104" -- 0CA4
           ,x"1304" -- 0CA6
           ,x"04c4" -- 0CA8
           ,x"05a0" -- 0CAA
           ,x"ec4c" -- 0CAC
           ,x"10f7" -- 0CAE
           ,x"05a0" -- 0CB0
           ,x"ec4e" -- 0CB2
           ,x"c0a0" -- 0CB4
           ,x"ec4e" -- 0CB6
           ,x"0a22" -- 0CB8
           ,x"0222" -- 0CBA
           ,x"ec62" -- 0CBC
           ,x"0642" -- 0CBE
           ,x"ccb0" -- 0CC0
           ,x"c4b0" -- 0CC2
           ,x"045c" -- 0CC4
           ,x"0000" -- 0CC6
           ,x"0a00" -- 0CC8
           ,x"0a9a" -- 0CCA
           ,x"0a66" -- 0CCC
           ,x"0a5e" -- 0CCE
           ,x"0aa0" -- 0CD0
           ,x"0ac8" -- 0CD2
           ,x"088e" -- 0CD4
           ,x"0905" -- 0CD6
           ,x"0a0a" -- 0CD8
           ,x"1408" -- 0CDA
           ,x"0013" -- 0CDC
           ,x"0a06" -- 0CDE
           ,x"0310" -- 0CE0
           ,x"0307" -- 0CE2
           ,x"0122" -- 0CE4
           ,x"5329" -- 0CE6
           ,x"aec4" -- 0CE8
           ,x"69af" -- 0CEA
           ,x"d267" -- 0CEC
           ,x"022c" -- 0CEE
           ,x"d770" -- 0CF0
           ,x"b353" -- 0CF2
           ,x"0322" -- 0CF4
           ,x"29ab" -- 0CF6
           ,x"cf6e" -- 0CF8
           ,x"66ac" -- 0CFA
           ,x"52af" -- 0CFC
           ,x"43ba" -- 0CFE
           ,x"4384" -- 0D00
           ,x"a1d4" -- 0D02
           ,x"61a5" -- 0D04
           ,x"4374" -- 0D06
           ,x"a956" -- 0D08
           ,x"7385" -- 0D0A
           ,x"ae44" -- 0D0C
           ,x"b155" -- 0D0E
           ,x"89a4" -- 0D10
           ,x"cc65" -- 0D12
           ,x"ae43" -- 0D14
           ,x"7456" -- 0D16
           ,x"8aa5" -- 0D18
           ,x"51a7" -- 0D1A
           ,x"5428" -- 0D1C
           ,x"452c" -- 0D1E
           ,x"4554" -- 0D20
           ,x"ad50" -- 0D22
           ,x"ae43" -- 0D24
           ,x"454f" -- 0D26
           ,x"af43" -- 0D28
           ,x"508c" -- 0D2A
           ,x"a4c3" -- 0D2C
           ,x"7229" -- 0D2E
           ,x"cd69" -- 0D30
           ,x"b2c5" -- 0D32
           ,x"78b3" -- 0D34
           ,x"54b7" -- 0D36
           ,x"5069" -- 0D38
           ,x"8daf" -- 0D3A
           ,x"5662" -- 0D3C
           ,x"b059" -- 0D3E
           ,x"738e" -- 0D40
           ,x"a547" -- 0D42
           ,x"af50" -- 0D44
           ,x"8fb2" -- 0D46
           ,x"4992" -- 0D48
           ,x"b3c5" -- 0D4A
           ,x"74b4" -- 0D4C
           ,x"d770" -- 0D4E
           ,x"1322" -- 0D50
           ,x"4f5a" -- 0D52
           ,x"a5d4" -- 0D54
           ,x"6fac" -- 0D56
           ,x"41af" -- 0D58
           ,x"4362" -- 0D5A
           ,x"b241" -- 0D5C
           ,x"434c" -- 0D5E
           ,x"b4c3" -- 0D60
           ,x"72d3" -- 0D62
           ,x"74d7" -- 0D64
           ,x"70b7" -- 0D66
           ,x"d062" -- 0D68
           ,x"ba43" -- 0D6A
           ,x"6294" -- 0D6C
           ,x"22a5" -- 0D6E
           ,x"d874" -- 0D70
           ,x"18af" -- 0D72
           ,x"5052" -- 0D74
           ,x"0000" -- 0D76
           ,x"a000" -- 0D78
           ,x"b000" -- 0D7A
           ,x"0745" -- 0D7C
           ,x"0227" -- 0D7E
           ,x"0247" -- 0D80
           ,x"000d" -- 0D82
           ,x"0445" -- 0D84
           ,x"0685" -- 0D86
           ,x"0405" -- 0D88
           ,x"000d" -- 0D8A
           ,x"8000" -- 0D8C
           ,x"9000" -- 0D8E
           ,x"0287" -- 0D90
           ,x"03a6" -- 0D92
           ,x"03c6" -- 0D94
           ,x"04c5" -- 0D96
           ,x"2002" -- 0D98
           ,x"2402" -- 0D9A
           ,x"000a" -- 0D9C
           ,x"0605" -- 0D9E
           ,x"0645" -- 0DA0
           ,x"3c08" -- 0DA2
           ,x"0185" -- 0DA4
           ,x"000c" -- 0DA6
           ,x"0006" -- 0DA8
           ,x"0346" -- 0DAA
           ,x"0585" -- 0DAC
           ,x"05c5" -- 0DAE
           ,x"0545" -- 0DB0
           ,x"1301" -- 0DB2
           ,x"1501" -- 0DB4
           ,x"1b01" -- 0DB6
           ,x"1401" -- 0DB8
           ,x"1a01" -- 0DBA
           ,x"1201" -- 0DBC
           ,x"1101" -- 0DBE
           ,x"1001" -- 0DC0
           ,x"1701" -- 0DC2
           ,x"1601" -- 0DC4
           ,x"1901" -- 0DC6
           ,x"1801" -- 0DC8
           ,x"1c01" -- 0DCA
           ,x"3003" -- 0DCC
           ,x"0207" -- 0DCE
           ,x"030a" -- 0DD0
           ,x"03e6" -- 0DD2
           ,x"008b" -- 0DD4
           ,x"009b" -- 0DD6
           ,x"02ea" -- 0DD8
           ,x"c000" -- 0DDA
           ,x"d000" -- 0DDC
           ,x"3808" -- 0DDE
           ,x"01c5" -- 0DE0
           ,x"0505" -- 0DE2
           ,x"1006" -- 0DE4
           ,x"0267" -- 0DE6
           ,x"0366" -- 0DE8
           ,x"0386" -- 0DEA
           ,x"6000" -- 0DEC
           ,x"7000" -- 0DEE
           ,x"1d09" -- 0DF0
           ,x"1e09" -- 0DF2
           ,x"0705" -- 0DF4
           ,x"0a04" -- 0DF6
           ,x"e000" -- 0DF8
           ,x"f000" -- 0DFA
           ,x"0804" -- 0DFC
           ,x"0b04" -- 0DFE
           ,x"0904" -- 0E00
           ,x"3403" -- 0E02
           ,x"02cb" -- 0E04
           ,x"02ab" -- 0E06
           ,x"06c5" -- 0E08
           ,x"4000" -- 0E0A
           ,x"5000" -- 0E0C
           ,x"1f09" -- 0E0E
           ,x"0006" -- 0E10
           ,x"0485" -- 0E12
           ,x"2c08" -- 0E14
           ,x"2802" -- 0E16
           ,x"0000" -- 0E18
           ,x"02e0" -- 0E1A
           ,x"ec00" -- 0E1C
           ,x"0203" -- 0E1E
           ,x"ec4c" -- 0E20
           ,x"0205" -- 0E22
           ,x"ed00" -- 0E24
           ,x"0206" -- 0E26
           ,x"effe" -- 0E28
           ,x"ccc5" -- 0E2A
           ,x"ccc6" -- 0E2C
           ,x"ccc5" -- 0E2E
           ,x"04c5" -- 0E30
           ,x"04d3" -- 0E32
           ,x"0209" -- 0E34
           ,x"ec2e" -- 0E36
           ,x"c820" -- 0E38
           ,x"ec44" -- 0E3A
           ,x"ec54" -- 0E3C
           ,x"020c" -- 0E3E
           ,x"0400" -- 0E40
           ,x"1d1f" -- 0E42
           ,x"3220" -- 0E44
           ,x"013b" -- 0E46
           ,x"1e0d" -- 0E48
           ,x"3320" -- 0E4A
           ,x"0096" -- 0E4C
           ,x"1d10" -- 0E4E
           ,x"020c" -- 0E50
           ,x"0000" -- 0E52
           ,x"1d0e" -- 0E54
           ,x"3220" -- 0E56
           ,x"013b" -- 0E58
           ,x"04c1" -- 0E5A
           ,x"04c2" -- 0E5C
           ,x"c660" -- 0E5E
           ,x"013e" -- 0E60
           ,x"2fa0" -- 0E62
           ,x"00e3" -- 0E64
           ,x"05e0" -- 0E66
           ,x"ec44" -- 0E68
           ,x"020c" -- 0E6A
           ,x"0000" -- 0E6C
           ,x"1f15" -- 0E6E
           ,x"1334" -- 0E70
           ,x"020c" -- 0E72
           ,x"0400" -- 0E74
           ,x"1f15" -- 0E76
           ,x"1303" -- 0E78
           ,x"c041" -- 0E7A
           ,x"162c" -- 0E7C
           ,x"10f5" -- 0E7E
           ,x"c660" -- 0E80
           ,x"0140" -- 0E82
           ,x"c082" -- 0E84
           ,x"1625" -- 0E86
           ,x"2f4a" -- 0E88
           ,x"028a" -- 0E8A
           ,x"0000" -- 0E8C
           ,x"13ed" -- 0E8E
           ,x"028a" -- 0E90
           ,x"7f00" -- 0E92
           ,x"13ea" -- 0E94
           ,x"028a" -- 0E96
           ,x"1000" -- 0E98
           ,x"160d" -- 0E9A
           ,x"2f4a" -- 0E9C
           ,x"028a" -- 0E9E
           ,x"0000" -- 0EA0
           ,x"13fc" -- 0EA2
           ,x"028a" -- 0EA4
           ,x"3700" -- 0EA6
           ,x"130e" -- 0EA8
           ,x"028a" -- 0EAA
           ,x"3c00" -- 0EAC
           ,x"16dd" -- 0EAE
           ,x"2f20" -- 0EB0
           ,x"013c" -- 0EB2
           ,x"10da" -- 0EB4
           ,x"028a" -- 0EB6
           ,x"1200" -- 0EB8
           ,x"1602" -- 0EBA
           ,x"0460" -- 0EBC
           ,x"1070" -- 0EBE
           ,x"028a" -- 0EC0
           ,x"1100" -- 0EC2
           ,x"1602" -- 0EC4
           ,x"0460" -- 0EC6
           ,x"0fa0" -- 0EC8
           ,x"c660" -- 0ECA
           ,x"013e" -- 0ECC
           ,x"2f0a" -- 0ECE
           ,x"10cc" -- 0ED0
           ,x"0460" -- 0ED2
           ,x"107c" -- 0ED4
           ,x"0460" -- 0ED6
           ,x"0fc8" -- 0ED8
           ,x"c660" -- 0EDA
           ,x"013e" -- 0EDC
           ,x"2f4a" -- 0EDE
           ,x"028a" -- 0EE0
           ,x"1a00" -- 0EE2
           ,x"1605" -- 0EE4
           ,x"c820" -- 0EE6
           ,x"ec54" -- 0EE8
           ,x"ec44" -- 0EEA
           ,x"0460" -- 0EEC
           ,x"0142" -- 0EEE
           ,x"028a" -- 0EF0
           ,x"0300" -- 0EF2
           ,x"1310" -- 0EF4
           ,x"028a" -- 0EF6
           ,x"1200" -- 0EF8
           ,x"13e0" -- 0EFA
           ,x"028a" -- 0EFC
           ,x"1400" -- 0EFE
           ,x"1602" -- 0F00
           ,x"0460" -- 0F02
           ,x"10fe" -- 0F04
           ,x"c041" -- 0F06
           ,x"16e6" -- 0F08
           ,x"c082" -- 0F0A
           ,x"16e2" -- 0F0C
           ,x"c660" -- 0F0E
           ,x"0140" -- 0F10
           ,x"2f0a" -- 0F12
           ,x"10aa" -- 0F14
           ,x"c660" -- 0F16
           ,x"013e" -- 0F18
           ,x"c820" -- 0F1A
           ,x"ec54" -- 0F1C
           ,x"ec44" -- 0F1E
           ,x"2fa0" -- 0F20
           ,x"00d8" -- 0F22
           ,x"2eca" -- 0F24
           ,x"2fa0" -- 0F26
           ,x"00de" -- 0F28
           ,x"06a0" -- 0F2A
           ,x"0f42" -- 0F2C
           ,x"5500" -- 0F2E
           ,x"0f7e" -- 0F30
           ,x"4400" -- 0F32
           ,x"0f94" -- 0F34
           ,x"5400" -- 0F36
           ,x"0f5a" -- 0F38
           ,x"5100" -- 0F3A
           ,x"0e5a" -- 0F3C
           ,x"0000" -- 0F3E
           ,x"05cb" -- 0F40
           ,x"c01b" -- 0F42
           ,x"1304" -- 0F44
           ,x"82bb" -- 0F46
           ,x"16fb" -- 0F48
           ,x"c2db" -- 0F4A
           ,x"045b" -- 0F4C
           ,x"2fa0" -- 0F4E
           ,x"00f5" -- 0F50
           ,x"10e1" -- 0F52
           ,x"2fa0" -- 0F54
           ,x"00ff" -- 0F56
           ,x"10de" -- 0F58
           ,x"2e4a" -- 0F5A
           ,x"0f16" -- 0F5C
           ,x"0f54" -- 0F5E
           ,x"0a2a" -- 0F60
           ,x"064a" -- 0F62
           ,x"12f7" -- 0F64
           ,x"028a" -- 0F66
           ,x"0023" -- 0F68
           ,x"14f4" -- 0F6A
           ,x"020c" -- 0F6C
           ,x"0400" -- 0F6E
           ,x"1d0b" -- 0F70
           ,x"1d0c" -- 0F72
           ,x"332a" -- 0F74
           ,x"0084" -- 0F76
           ,x"1e0b" -- 0F78
           ,x"1e0c" -- 0F7A
           ,x"10cc" -- 0F7C
           ,x"2e4a" -- 0F7E
           ,x"0f88" -- 0F80
           ,x"0f54" -- 0F82
           ,x"c80a" -- 0F84
           ,x"ec50" -- 0F86
           ,x"2e4a" -- 0F88
           ,x"0f16" -- 0F8A
           ,x"0f54" -- 0F8C
           ,x"c80a" -- 0F8E
           ,x"ec4e" -- 0F90
           ,x"10c1" -- 0F92
           ,x"2e4a" -- 0F94
           ,x"0f16" -- 0F96
           ,x"0f54" -- 0F98
           ,x"c80a" -- 0F9A
           ,x"ec4c" -- 0F9C
           ,x"10bb" -- 0F9E
           ,x"0701" -- 0FA0
           ,x"c1e0" -- 0FA2
           ,x"ec52" -- 0FA4
           ,x"112d" -- 0FA6
           ,x"1533" -- 0FA8
           ,x"c1e0" -- 0FAA
           ,x"ec50" -- 0FAC
           ,x"8807" -- 0FAE
           ,x"ec4e" -- 0FB0
           ,x"1b37" -- 0FB2
           ,x"c660" -- 0FB4
           ,x"0140" -- 0FB6
           ,x"04c5" -- 0FB8
           ,x"04c3" -- 0FBA
           ,x"2fa0" -- 0FBC
           ,x"0137" -- 0FBE
           ,x"c287" -- 0FC0
           ,x"06a0" -- 0FC2
           ,x"1042" -- 0FC4
           ,x"3900" -- 0FC6
           ,x"c297" -- 0FC8
           ,x"06a0" -- 0FCA
           ,x"1042" -- 0FCC
           ,x"4200" -- 0FCE
           ,x"8807" -- 0FD0
           ,x"ec4e" -- 0FD2
           ,x"1a03" -- 0FD4
           ,x"0720" -- 0FD6
           ,x"ec52" -- 0FD8
           ,x"1004" -- 0FDA
           ,x"05c7" -- 0FDC
           ,x"0283" -- 0FDE
           ,x"003c" -- 0FE0
           ,x"111d" -- 0FE2
           ,x"0225" -- 0FE4
           ,x"0037" -- 0FE6
           ,x"c285" -- 0FE8
           ,x"050a" -- 0FEA
           ,x"06a0" -- 0FEC
           ,x"1042" -- 0FEE
           ,x"3700" -- 0FF0
           ,x"c807" -- 0FF2
           ,x"ec50" -- 0FF4
           ,x"2fa0" -- 0FF6
           ,x"0128" -- 0FF8
           ,x"c160" -- 0FFA
           ,x"ec54" -- 0FFC
           ,x"110e" -- 0FFE
           ,x"10cf" -- 1000
           ,x"2fa0" -- 1002
           ,x"0137" -- 1004
           ,x"2fa0" -- 1006
           ,x"00e0" -- 1008
           ,x"05e0" -- 100A
           ,x"ec52" -- 100C
           ,x"10f5" -- 100E
           ,x"2fa0" -- 1010
           ,x"0137" -- 1012
           ,x"2fa0" -- 1014
           ,x"0131" -- 1016
           ,x"04e0" -- 1018
           ,x"ec52" -- 101A
           ,x"04c1" -- 101C
           ,x"0460" -- 101E
           ,x"0e6a" -- 1020
           ,x"2fa0" -- 1022
           ,x"0137" -- 1024
           ,x"2fa0" -- 1026
           ,x"0131" -- 1028
           ,x"c660" -- 102A
           ,x"013e" -- 102C
           ,x"c820" -- 102E
           ,x"ec54" -- 1030
           ,x"ec44" -- 1032
           ,x"2fa0" -- 1034
           ,x"011f" -- 1036
           ,x"05e0" -- 1038
           ,x"ec44" -- 103A
           ,x"0720" -- 103C
           ,x"ec4c" -- 103E
           ,x"10eb" -- 1040
           ,x"c03b" -- 1042
           ,x"2f00" -- 1044
           ,x"0980" -- 1046
           ,x"a140" -- 1048
           ,x"2e8a" -- 104A
           ,x"0223" -- 104C
           ,x"0005" -- 104E
           ,x"0200" -- 1050
           ,x"0004" -- 1052
           ,x"0b4a" -- 1054
           ,x"c18a" -- 1056
           ,x"09c6" -- 1058
           ,x"a146" -- 105A
           ,x"0225" -- 105C
           ,x"0030" -- 105E
           ,x"0286" -- 1060
           ,x"000a" -- 1062
           ,x"1a02" -- 1064
           ,x"0225" -- 1066
           ,x"0007" -- 1068
           ,x"0600" -- 106A
           ,x"16f3" -- 106C
           ,x"045b" -- 106E
           ,x"0702" -- 1070
           ,x"c660" -- 1072
           ,x"0140" -- 1074
           ,x"c020" -- 1076
           ,x"ec4c" -- 1078
           ,x"04c7" -- 107A
           ,x"2f46" -- 107C
           ,x"0286" -- 107E
           ,x"1400" -- 1080
           ,x"133d" -- 1082
           ,x"c220" -- 1084
           ,x"ec52" -- 1086
           ,x"1657" -- 1088
           ,x"0286" -- 108A
           ,x"2000" -- 108C
           ,x"11f6" -- 108E
           ,x"0286" -- 1090
           ,x"5f00" -- 1092
           ,x"15f3" -- 1094
           ,x"0705" -- 1096
           ,x"04ca" -- 1098
           ,x"06a0" -- 109A
           ,x"073a" -- 109C
           ,x"100b" -- 109E
           ,x"d22a" -- 10A0
           ,x"1152" -- 10A2
           ,x"1332" -- 10A4
           ,x"06a0" -- 10A6
           ,x"0722" -- 10A8
           ,x"100e" -- 10AA
           ,x"0205" -- 10AC
           ,x"0008" -- 10AE
           ,x"0878" -- 10B0
           ,x"0468" -- 10B2
           ,x"10b2" -- 10B4
           ,x"0286" -- 10B6
           ,x"0047" -- 10B8
           ,x"1106" -- 10BA
           ,x"0286" -- 10BC
           ,x"004a" -- 10BE
           ,x"1522" -- 10C0
           ,x"0226" -- 10C2
           ,x"ffc9" -- 10C4
           ,x"10ec" -- 10C6
           ,x"0286" -- 10C8
           ,x"003a" -- 10CA
           ,x"161c" -- 10CC
           ,x"103e" -- 10CE
           ,x"020c" -- 10D0
           ,x"0400" -- 10D2
           ,x"04c5" -- 10D4
           ,x"1f0f" -- 10D6
           ,x"16fd" -- 10D8
           ,x"0605" -- 10DA
           ,x"16fc" -- 10DC
           ,x"c660" -- 10DE
           ,x"013e" -- 10E0
           ,x"c820" -- 10E2
           ,x"ec54" -- 10E4
           ,x"ec44" -- 10E6
           ,x"0720" -- 10E8
           ,x"ec4c" -- 10EA
           ,x"c000" -- 10EC
           ,x"1303" -- 10EE
           ,x"2fa0" -- 10F0
           ,x"010a" -- 10F2
           ,x"1002" -- 10F4
           ,x"2fa0" -- 10F6
           ,x"0115" -- 10F8
           ,x"05e0" -- 10FA
           ,x"ec44" -- 10FC
           ,x"04c2" -- 10FE
           ,x"04e0" -- 1100
           ,x"ec52" -- 1102
           ,x"1021" -- 1104
           ,x"04c0" -- 1106
           ,x"10e3" -- 1108
           ,x"2f46" -- 110A
           ,x"9806" -- 110C
           ,x"00f2" -- 110E
           ,x"16fc" -- 1110
           ,x"04c7" -- 1112
           ,x"1019" -- 1114
           ,x"a1ca" -- 1116
           ,x"1317" -- 1118
           ,x"0700" -- 111A
           ,x"10d9" -- 111C
           ,x"a280" -- 111E
           ,x"c0ca" -- 1120
           ,x"1012" -- 1122
           ,x"a280" -- 1124
           ,x"ccca" -- 1126
           ,x"100f" -- 1128
           ,x"0645" -- 112A
           ,x"2f46" -- 112C
           ,x"0986" -- 112E
           ,x"13fd" -- 1130
           ,x"a1c6" -- 1132
           ,x"0605" -- 1134
           ,x"16fa" -- 1136
           ,x"1007" -- 1138
           ,x"a280" -- 113A
           ,x"c80a" -- 113C
           ,x"ec1c" -- 113E
           ,x"1003" -- 1140
           ,x"024a" -- 1142
           ,x"fffe" -- 1144
           ,x"c00a" -- 1146
           ,x"0460" -- 1148
           ,x"0e6a" -- 114A
           ,x"0720" -- 114C
           ,x"ec52" -- 114E
           ,x"10fb" -- 1150
           ,x"3d45" -- 1152
           ,x"443c" -- 1154
           ,x"3c3c" -- 1156
           ,x"3c32" -- 1158
           ,x"e437" -- 115A
           ,x"363a" -- 115C
           ,x"3948" -- 115E
           ,x"2a00" -- 1160
           ,x"3c3c" -- 1162
           ,x"3d8b" -- 1164
           ,x"c141" -- 1166
           ,x"0208" -- 1168
           ,x"12d8" -- 116A
           ,x"0209" -- 116C
           ,x"12ba" -- 116E
           ,x"0207" -- 1170
           ,x"12a6" -- 1172
           ,x"2fa0" -- 1174
           ,x"00f2" -- 1176
           ,x"0206" -- 1178
           ,x"202c" -- 117A
           ,x"c050" -- 117C
           ,x"2e80" -- 117E
           ,x"2f06" -- 1180
           ,x"2e81" -- 1182
           ,x"2f06" -- 1184
           ,x"04c3" -- 1186
           ,x"c050" -- 1188
           ,x"0241" -- 118A
           ,x"fff0" -- 118C
           ,x"c2a3" -- 118E
           ,x"13b4" -- 1190
           ,x"c08a" -- 1192
           ,x"1329" -- 1194
           ,x"024a" -- 1196
           ,x"fff0" -- 1198
           ,x"8281" -- 119A
           ,x"1402" -- 119C
           ,x"0643" -- 119E
           ,x"10f6" -- 11A0
           ,x"c050" -- 11A2
           ,x"0a13" -- 11A4
           ,x"0223" -- 11A6
           ,x"14d6" -- 11A8
           ,x"604a" -- 11AA
           ,x"0242" -- 11AC
           ,x"000f" -- 11AE
           ,x"d0a2" -- 11B0
           ,x"11ba" -- 11B2
           ,x"0972" -- 11B4
           ,x"0462" -- 11B6
           ,x"11ba" -- 11B8
           ,x"060c" -- 11BA
           ,x"061f" -- 11BC
           ,x"232b" -- 11BE
           ,x"3337" -- 11C0
           ,x"063f" -- 11C2
           ,x"4145" -- 11C4
           ,x"0697" -- 11C6
           ,x"0698" -- 11C8
           ,x"2f06" -- 11CA
           ,x"0961" -- 11CC
           ,x"0698" -- 11CE
           ,x"103d" -- 11D0
           ,x"c041" -- 11D2
           ,x"1603" -- 11D4
           ,x"0203" -- 11D6
           ,x"14da" -- 11D8
           ,x"1024" -- 11DA
           ,x"06c1" -- 11DC
           ,x"0871" -- 11DE
           ,x"05c1" -- 11E0
           ,x"a040" -- 11E2
           ,x"0697" -- 11E4
           ,x"1004" -- 11E6
           ,x"c050" -- 11E8
           ,x"0203" -- 11EA
           ,x"14de" -- 11EC
           ,x"0697" -- 11EE
           ,x"2f20" -- 11F0
           ,x"14f5" -- 11F2
           ,x"2e81" -- 11F4
           ,x"102a" -- 11F6
           ,x"0697" -- 11F8
           ,x"0698" -- 11FA
           ,x"c209" -- 11FC
           ,x"10e5" -- 11FE
           ,x"d041" -- 1200
           ,x"16f2" -- 1202
           ,x"0b41" -- 1204
           ,x"d081" -- 1206
           ,x"0a61" -- 1208
           ,x"09c2" -- 120A
           ,x"a042" -- 120C
           ,x"10f4" -- 120E
           ,x"8810" -- 1210
           ,x"1320" -- 1212
           ,x"1603" -- 1214
           ,x"0203" -- 1216
           ,x"14ee" -- 1218
           ,x"1004" -- 121A
           ,x"0697" -- 121C
           ,x"10d7" -- 121E
           ,x"c041" -- 1220
           ,x"16e2" -- 1222
           ,x"0697" -- 1224
           ,x"1012" -- 1226
           ,x"0ac1" -- 1228
           ,x"18de" -- 122A
           ,x"09c1" -- 122C
           ,x"0697" -- 122E
           ,x"0698" -- 1230
           ,x"2f06" -- 1232
           ,x"c070" -- 1234
           ,x"10dc" -- 1236
           ,x"0697" -- 1238
           ,x"1019" -- 123A
           ,x"c041" -- 123C
           ,x"16d4" -- 123E
           ,x"0697" -- 1240
           ,x"10f8" -- 1242
           ,x"0ac1" -- 1244
           ,x"18d0" -- 1246
           ,x"09c1" -- 1248
           ,x"10e2" -- 124A
           ,x"c145" -- 124C
           ,x"1603" -- 124E
           ,x"c740" -- 1250
           ,x"0460" -- 1252
           ,x"0142" -- 1254
           ,x"c320" -- 1256
           ,x"013e" -- 1258
           ,x"1f15" -- 125A
           ,x"1604" -- 125C
           ,x"2f42" -- 125E
           ,x"0282" -- 1260
           ,x"2f00" -- 1262
           ,x"13f5" -- 1264
           ,x"8140" -- 1266
           ,x"1bf3" -- 1268
           ,x"0460" -- 126A
           ,x"1168" -- 126C
           ,x"0203" -- 126E
           ,x"2d31" -- 1270
           ,x"06c1" -- 1272
           ,x"0881" -- 1274
           ,x"1315" -- 1276
           ,x"1502" -- 1278
           ,x"2f03" -- 127A
           ,x"0501" -- 127C
           ,x"0281" -- 127E
           ,x"0064" -- 1280
           ,x"1104" -- 1282
           ,x"0a83" -- 1284
           ,x"2f03" -- 1286
           ,x"0221" -- 1288
           ,x"ff9c" -- 128A
           ,x"0204" -- 128C
           ,x"000a" -- 128E
           ,x"c081" -- 1290
           ,x"04c1" -- 1292
           ,x"3c44" -- 1294
           ,x"0a83" -- 1296
           ,x"1302" -- 1298
           ,x"c041" -- 129A
           ,x"1301" -- 129C
           ,x"0699" -- 129E
           ,x"c042" -- 12A0
           ,x"0699" -- 12A2
           ,x"10d3" -- 12A4
           ,x"0202" -- 12A6
           ,x"0004" -- 12A8
           ,x"2f13" -- 12AA
           ,x"0583" -- 12AC
           ,x"0602" -- 12AE
           ,x"16fc" -- 12B0
           ,x"2f06" -- 12B2
           ,x"06c6" -- 12B4
           ,x"05c0" -- 12B6
           ,x"045b" -- 12B8
           ,x"c0c1" -- 12BA
           ,x"0ac3" -- 12BC
           ,x"0943" -- 12BE
           ,x"0283" -- 12C0
           ,x"0900" -- 12C2
           ,x"1203" -- 12C4
           ,x"06c3" -- 12C6
           ,x"0223" -- 12C8
           ,x"0126" -- 12CA
           ,x"0223" -- 12CC
           ,x"3000" -- 12CE
           ,x"2f03" -- 12D0
           ,x"0a83" -- 12D2
           ,x"16fd" -- 12D4
           ,x"045b" -- 12D6
           ,x"0204" -- 12D8
           ,x"2a52" -- 12DA
           ,x"c081" -- 12DC
           ,x"0aa2" -- 12DE
           ,x"09e2" -- 12E0
           ,x"1603" -- 12E2
           ,x"06c4" -- 12E4
           ,x"2f04" -- 12E6
           ,x"10e8" -- 12E8
           ,x"0602" -- 12EA
           ,x"1602" -- 12EC
           ,x"2f04" -- 12EE
           ,x"10f9" -- 12F0
           ,x"0602" -- 12F2
           ,x"1610" -- 12F4
           ,x"2fa0" -- 12F6
           ,x"14f4" -- 12F8
           ,x"2eb0" -- 12FA
           ,x"c081" -- 12FC
           ,x"0ac2" -- 12FE
           ,x"13ea" -- 1300
           ,x"0202" -- 1302
           ,x"2829" -- 1304
           ,x"2f02" -- 1306
           ,x"06c4" -- 1308
           ,x"2f04" -- 130A
           ,x"c30b" -- 130C
           ,x"0699" -- 130E
           ,x"06c2" -- 1310
           ,x"2f02" -- 1312
           ,x"045c" -- 1314
           ,x"2fa0" -- 1316
           ,x"14f7" -- 1318
           ,x"0202" -- 131A
           ,x"002b" -- 131C
           ,x"10f6" -- 131E
           ,x"045b" -- 1320
           ,x"0000" -- 1322
           ,x"008b" -- 1324
           ,x"009b" -- 1326
           ,x"0185" -- 1328
           ,x"01c5" -- 132A
           ,x"0207" -- 132C
           ,x"0227" -- 132E
           ,x"0247" -- 1330
           ,x"0267" -- 1332
           ,x"0287" -- 1334
           ,x"02ab" -- 1336
           ,x"02cb" -- 1338
           ,x"02ea" -- 133A
           ,x"030a" -- 133C
           ,x"0346" -- 133E
           ,x"0366" -- 1340
           ,x"0386" -- 1342
           ,x"03a6" -- 1344
           ,x"03c6" -- 1346
           ,x"03e6" -- 1348
           ,x"0405" -- 134A
           ,x"0445" -- 134C
           ,x"0485" -- 134E
           ,x"04c5" -- 1350
           ,x"0505" -- 1352
           ,x"0545" -- 1354
           ,x"0585" -- 1356
           ,x"05c5" -- 1358
           ,x"0605" -- 135A
           ,x"0645" -- 135C
           ,x"0685" -- 135E
           ,x"06c5" -- 1360
           ,x"0705" -- 1362
           ,x"0745" -- 1364
           ,x"0804" -- 1366
           ,x"0904" -- 1368
           ,x"0a04" -- 136A
           ,x"0b04" -- 136C
           ,x"1001" -- 136E
           ,x"1101" -- 1370
           ,x"1201" -- 1372
           ,x"1301" -- 1374
           ,x"1401" -- 1376
           ,x"1501" -- 1378
           ,x"1601" -- 137A
           ,x"1701" -- 137C
           ,x"1801" -- 137E
           ,x"1901" -- 1380
           ,x"1a01" -- 1382
           ,x"1b01" -- 1384
           ,x"1c01" -- 1386
           ,x"1d09" -- 1388
           ,x"1e09" -- 138A
           ,x"1f09" -- 138C
           ,x"2002" -- 138E
           ,x"2402" -- 1390
           ,x"2802" -- 1392
           ,x"2c03" -- 1394
           ,x"3003" -- 1396
           ,x"3403" -- 1398
           ,x"3808" -- 139A
           ,x"3c08" -- 139C
           ,x"4000" -- 139E
           ,x"5000" -- 13A0
           ,x"6000" -- 13A2
           ,x"7000" -- 13A4
           ,x"8000" -- 13A6
           ,x"9000" -- 13A8
           ,x"a000" -- 13AA
           ,x"b000" -- 13AC
           ,x"c000" -- 13AE
           ,x"d000" -- 13B0
           ,x"e000" -- 13B2
           ,x"f000" -- 13B4
           ,x"4c53" -- 13B6
           ,x"5420" -- 13B8
           ,x"4c57" -- 13BA
           ,x"5020" -- 13BC
           ,x"4449" -- 13BE
           ,x"5653" -- 13C0
           ,x"4d50" -- 13C2
           ,x"5953" -- 13C4
           ,x"4c49" -- 13C6
           ,x"2020" -- 13C8
           ,x"4149" -- 13CA
           ,x"2020" -- 13CC
           ,x"414e" -- 13CE
           ,x"4449" -- 13D0
           ,x"4f52" -- 13D2
           ,x"4920" -- 13D4
           ,x"4349" -- 13D6
           ,x"2020" -- 13D8
           ,x"5354" -- 13DA
           ,x"5750" -- 13DC
           ,x"5354" -- 13DE
           ,x"5354" -- 13E0
           ,x"4c57" -- 13E2
           ,x"5049" -- 13E4
           ,x"4c49" -- 13E6
           ,x"4d49" -- 13E8
           ,x"4944" -- 13EA
           ,x"4c45" -- 13EC
           ,x"5253" -- 13EE
           ,x"4554" -- 13F0
           ,x"5254" -- 13F2
           ,x"5750" -- 13F4
           ,x"434b" -- 13F6
           ,x"4f4e" -- 13F8
           ,x"434b" -- 13FA
           ,x"4f46" -- 13FC
           ,x"4c52" -- 13FE
           ,x"4558" -- 1400
           ,x"424c" -- 1402
           ,x"5750" -- 1404
           ,x"4220" -- 1406
           ,x"2020" -- 1408
           ,x"5820" -- 140A
           ,x"2020" -- 140C
           ,x"434c" -- 140E
           ,x"5220" -- 1410
           ,x"4e45" -- 1412
           ,x"4720" -- 1414
           ,x"494e" -- 1416
           ,x"5620" -- 1418
           ,x"494e" -- 141A
           ,x"4320" -- 141C
           ,x"494e" -- 141E
           ,x"4354" -- 1420
           ,x"4445" -- 1422
           ,x"4320" -- 1424
           ,x"4445" -- 1426
           ,x"4354" -- 1428
           ,x"424c" -- 142A
           ,x"2020" -- 142C
           ,x"5357" -- 142E
           ,x"5042" -- 1430
           ,x"5345" -- 1432
           ,x"544f" -- 1434
           ,x"4142" -- 1436
           ,x"5320" -- 1438
           ,x"5352" -- 143A
           ,x"4120" -- 143C
           ,x"5352" -- 143E
           ,x"4c20" -- 1440
           ,x"534c" -- 1442
           ,x"4120" -- 1444
           ,x"5352" -- 1446
           ,x"4320" -- 1448
           ,x"4a4d" -- 144A
           ,x"5020" -- 144C
           ,x"4a4c" -- 144E
           ,x"5420" -- 1450
           ,x"4a4c" -- 1452
           ,x"4520" -- 1454
           ,x"4a45" -- 1456
           ,x"5120" -- 1458
           ,x"4a48" -- 145A
           ,x"4520" -- 145C
           ,x"4a47" -- 145E
           ,x"5420" -- 1460
           ,x"4a4e" -- 1462
           ,x"4520" -- 1464
           ,x"4a4e" -- 1466
           ,x"4320" -- 1468
           ,x"4a4f" -- 146A
           ,x"4320" -- 146C
           ,x"4a4e" -- 146E
           ,x"4f20" -- 1470
           ,x"4a4c" -- 1472
           ,x"2020" -- 1474
           ,x"4a48" -- 1476
           ,x"2020" -- 1478
           ,x"4a4f" -- 147A
           ,x"5020" -- 147C
           ,x"5342" -- 147E
           ,x"4f20" -- 1480
           ,x"5342" -- 1482
           ,x"5a20" -- 1484
           ,x"5442" -- 1486
           ,x"2020" -- 1488
           ,x"434f" -- 148A
           ,x"4320" -- 148C
           ,x"435a" -- 148E
           ,x"4320" -- 1490
           ,x"584f" -- 1492
           ,x"5220" -- 1494
           ,x"584f" -- 1496
           ,x"5020" -- 1498
           ,x"4c44" -- 149A
           ,x"4352" -- 149C
           ,x"5354" -- 149E
           ,x"4352" -- 14A0
           ,x"4d50" -- 14A2
           ,x"5920" -- 14A4
           ,x"4449" -- 14A6
           ,x"5620" -- 14A8
           ,x"535a" -- 14AA
           ,x"4320" -- 14AC
           ,x"535a" -- 14AE
           ,x"4342" -- 14B0
           ,x"5320" -- 14B2
           ,x"2020" -- 14B4
           ,x"5342" -- 14B6
           ,x"2020" -- 14B8
           ,x"4320" -- 14BA
           ,x"2020" -- 14BC
           ,x"4342" -- 14BE
           ,x"2020" -- 14C0
           ,x"4120" -- 14C2
           ,x"2020" -- 14C4
           ,x"4142" -- 14C6
           ,x"2020" -- 14C8
           ,x"4d4f" -- 14CA
           ,x"5620" -- 14CC
           ,x"4d4f" -- 14CE
           ,x"5642" -- 14D0
           ,x"534f" -- 14D2
           ,x"4320" -- 14D4
           ,x"534f" -- 14D6
           ,x"4342" -- 14D8
           ,x"4e4f" -- 14DA
           ,x"5020" -- 14DC
           ,x"4441" -- 14DE
           ,x"5441" -- 14E0
           ,x"5445" -- 14E2
           ,x"5854" -- 14E4
           ,x"414f" -- 14E6
           ,x"5247" -- 14E8
           ,x"454e" -- 14EA
           ,x"4420" -- 14EC
           ,x"5254" -- 14EE
           ,x"2020" -- 14F0
           ,x"0000" -- 14F2
           ,x"403e" -- 14F4
           ,x"002a" -- 14F6
           ,x"5200" -- 14F8
           ,x"ffff" -- 14FA
           ,x"ffff" -- 14FC
           ,x"ffff" -- 14FE
           ,x"2fa0" -- 1500
           ,x"1530" -- 1502
           ,x"2f41" -- 1504
           ,x"0281" -- 1506
           ,x"3100" -- 1508
           ,x"1604" -- 150A
           ,x"2fa0" -- 150C
           ,x"00ad" -- 150E
           ,x"0460" -- 1510
           ,x"0142" -- 1512
           ,x"0281" -- 1514
           ,x"3200" -- 1516
           ,x"16f5" -- 1518
           ,x"0201" -- 151A
           ,x"1600" -- 151C
           ,x"0202" -- 151E
           ,x"8000" -- 1520
           ,x"0203" -- 1522
           ,x"5eba" -- 1524
           ,x"ccb1" -- 1526
           ,x"0643" -- 1528
           ,x"16fd" -- 152A
           ,x"0460" -- 152C
           ,x"8036" -- 152E
           ,x"0d0a" -- 1530
           ,x"544d" -- 1532
           ,x"5320" -- 1534
           ,x"3939" -- 1536
           ,x"3935" -- 1538
           ,x"2042" -- 153A
           ,x"5245" -- 153C
           ,x"4144" -- 153E
           ,x"424f" -- 1540
           ,x"4152" -- 1542
           ,x"4420" -- 1544
           ,x"5359" -- 1546
           ,x"5354" -- 1548
           ,x"454d" -- 154A
           ,x"0d0a" -- 154C
           ,x"4259" -- 154E
           ,x"2053" -- 1550
           ,x"5455" -- 1552
           ,x"4152" -- 1554
           ,x"5420" -- 1556
           ,x"434f" -- 1558
           ,x"4e4e" -- 155A
           ,x"4552" -- 155C
           ,x"0d0a" -- 155E
           ,x"0d0a" -- 1560
           ,x"5052" -- 1562
           ,x"4553" -- 1564
           ,x"5320" -- 1566
           ,x"3120" -- 1568
           ,x"464f" -- 156A
           ,x"5220" -- 156C
           ,x"4556" -- 156E
           ,x"4d42" -- 1570
           ,x"5547" -- 1572
           ,x"204d" -- 1574
           ,x"4f4e" -- 1576
           ,x"4954" -- 1578
           ,x"4f52" -- 157A
           ,x"0d0a" -- 157C
           ,x"5052" -- 157E
           ,x"4553" -- 1580
           ,x"5320" -- 1582
           ,x"3220" -- 1584
           ,x"464f" -- 1586
           ,x"5220" -- 1588
           ,x"434f" -- 158A
           ,x"5254" -- 158C
           ,x"4558" -- 158E
           ,x"2042" -- 1590
           ,x"4153" -- 1592
           ,x"4943" -- 1594
           ,x"0d0a" -- 1596
           ,x"0000" -- 1598
           ,x"ffff" -- 159A
           ,x"ffff" -- 159C
           ,x"ffff" -- 159E
           ,x"ffff" -- 15A0
           ,x"ffff" -- 15A2
           ,x"ffff" -- 15A4
           ,x"ffff" -- 15A6
           ,x"ffff" -- 15A8
           ,x"ffff" -- 15AA
           ,x"ffff" -- 15AC
           ,x"ffff" -- 15AE
           ,x"ffff" -- 15B0
           ,x"ffff" -- 15B2
           ,x"ffff" -- 15B4
           ,x"ffff" -- 15B6
           ,x"ffff" -- 15B8
           ,x"ffff" -- 15BA
           ,x"ffff" -- 15BC
           ,x"ffff" -- 15BE
           ,x"ffff" -- 15C0
           ,x"ffff" -- 15C2
           ,x"ffff" -- 15C4
           ,x"ffff" -- 15C6
           ,x"ffff" -- 15C8
           ,x"ffff" -- 15CA
           ,x"ffff" -- 15CC
           ,x"ffff" -- 15CE
           ,x"ffff" -- 15D0
           ,x"ffff" -- 15D2
           ,x"ffff" -- 15D4
           ,x"ffff" -- 15D6
           ,x"ffff" -- 15D8
           ,x"ffff" -- 15DA
           ,x"ffff" -- 15DC
           ,x"ffff" -- 15DE
           ,x"ffff" -- 15E0
           ,x"ffff" -- 15E2
           ,x"ffff" -- 15E4
           ,x"ffff" -- 15E6
           ,x"ffff" -- 15E8
           ,x"ffff" -- 15EA
           ,x"ffff" -- 15EC
           ,x"ffff" -- 15EE
           ,x"ffff" -- 15F0
           ,x"ffff" -- 15F2
           ,x"ffff" -- 15F4
           ,x"ffff" -- 15F6
           ,x"ffff" -- 15F8
           ,x"ffff" -- 15FA
           ,x"ffff" -- 15FC
           ,x"ffff" -- 15FE
           ,x"ed1e" -- 1600
           ,x"ed24" -- 1602
           ,x"ed2e" -- 1604
           ,x"ed00" -- 1606
           ,x"edee" -- 1608
           ,x"edf8" -- 160A
           ,x"b4b2" -- 160C
           ,x"ed3a" -- 160E
           ,x"803a" -- 1610
           ,x"ef60" -- 1612
           ,x"ef68" -- 1614
           ,x"ef88" -- 1616
           ,x"efa8" -- 1618
           ,x"efaa" -- 161A
           ,x"efac" -- 161C
           ,x"efae" -- 161E
           ,x"efb0" -- 1620
           ,x"efb2" -- 1622
           ,x"efb4" -- 1624
           ,x"efbe" -- 1626
           ,x"efc4" -- 1628
           ,x"efc6" -- 162A
           ,x"8040" -- 162C
           ,x"8042" -- 162E
           ,x"0000" -- 1630
           ,x"0000" -- 1632
           ,x"0000" -- 1634
           ,x"0460" -- 1636
           ,x"cc94" -- 1638
           ,x"0000" -- 163A
           ,x"0000" -- 163C
           ,x"0000" -- 163E
           ,x"0000" -- 1640
           ,x"0000" -- 1642
           ,x"0000" -- 1644
           ,x"0000" -- 1646
           ,x"0000" -- 1648
           ,x"0000" -- 164A
           ,x"0000" -- 164C
           ,x"ffff" -- 164E
           ,x"ffff" -- 1650
           ,x"8142" -- 1652
           ,x"ffff" -- 1654
           ,x"ffff" -- 1656
           ,x"ffff" -- 1658
           ,x"ffff" -- 165A
           ,x"ffff" -- 165C
           ,x"ed3e" -- 165E
           ,x"ffff" -- 1660
           ,x"8084" -- 1662
           ,x"851a" -- 1664
           ,x"d050" -- 1666
           ,x"0000" -- 1668
           ,x"0000" -- 166A
           ,x"0000" -- 166C
           ,x"0000" -- 166E
           ,x"0000" -- 1670
           ,x"0000" -- 1672
           ,x"0000" -- 1674
           ,x"0000" -- 1676
           ,x"0000" -- 1678
           ,x"0000" -- 167A
           ,x"0000" -- 167C
           ,x"0000" -- 167E
           ,x"0000" -- 1680
           ,x"0000" -- 1682
           ,x"0001" -- 1684
           ,x"0203" -- 1686
           ,x"0405" -- 1688
           ,x"0607" -- 168A
           ,x"0809" -- 168C
           ,x"0a0b" -- 168E
           ,x"0c0d" -- 1690
           ,x"0e0f" -- 1692
           ,x"c820" -- 1694
           ,x"b920" -- 1696
           ,x"8044" -- 1698
           ,x"05a0" -- 169A
           ,x"8044" -- 169C
           ,x"d820" -- 169E
           ,x"c84c" -- 16A0
           ,x"ed91" -- 16A2
           ,x"0420" -- 16A4
           ,x"819c" -- 16A6
           ,x"04e0" -- 16A8
           ,x"8030" -- 16AA
           ,x"04e0" -- 16AC
           ,x"8032" -- 16AE
           ,x"04e0" -- 16B0
           ,x"ed36" -- 16B2
           ,x"045b" -- 16B4
           ,x"0420" -- 16B6
           ,x"8d70" -- 16B8
           ,x"0032" -- 16BA
           ,x"4300" -- 16BC
           ,x"0420" -- 16BE
           ,x"8d70" -- 16C0
           ,x"0031" -- 16C2
           ,x"c060" -- 16C4
           ,x"ed10" -- 16C6
           ,x"06a0" -- 16C8
           ,x"b52a" -- 16CA
           ,x"100c" -- 16CC
           ,x"c820" -- 16CE
           ,x"801c" -- 16D0
           ,x"ef9e" -- 16D2
           ,x"0420" -- 16D4
           ,x"b558" -- 16D6
           ,x"8802" -- 16D8
           ,x"ed04" -- 16DA
           ,x"14f0" -- 16DC
           ,x"8802" -- 16DE
           ,x"8048" -- 16E0
           ,x"1aed" -- 16E2
           ,x"c042" -- 16E4
           ,x"c801" -- 16E6
           ,x"ed10" -- 16E8
           ,x"c801" -- 16EA
           ,x"ed0e" -- 16EC
           ,x"020b" -- 16EE
           ,x"814a" -- 16F0
           ,x"c060" -- 16F2
           ,x"ed0e" -- 16F4
           ,x"c801" -- 16F6
           ,x"edd2" -- 16F8
           ,x"04f1" -- 16FA
           ,x"c801" -- 16FC
           ,x"edd4" -- 16FE
           ,x"c0c1" -- 1700
           ,x"0223" -- 1702
           ,x"0008" -- 1704
           ,x"c803" -- 1706
           ,x"edd6" -- 1708
           ,x"0223" -- 170A
           ,x"0008" -- 170C
           ,x"c803" -- 170E
           ,x"edd8" -- 1710
           ,x"0460" -- 1712
           ,x"ae9a" -- 1714
           ,x"0201" -- 1716
           ,x"c8b1" -- 1718
           ,x"04e0" -- 171A
           ,x"ede0" -- 171C
           ,x"04e0" -- 171E
           ,x"ed30" -- 1720
           ,x"1002" -- 1722
           ,x"0201" -- 1724
           ,x"c8b9" -- 1726
           ,x"04e0" -- 1728
           ,x"ede4" -- 172A
           ,x"04e0" -- 172C
           ,x"8046" -- 172E
           ,x"04e0" -- 1730
           ,x"edf0" -- 1732
           ,x"0420" -- 1734
           ,x"8178" -- 1736
           ,x"06a0" -- 1738
           ,x"c02c" -- 173A
           ,x"06a0" -- 173C
           ,x"a374" -- 173E
           ,x"10f1" -- 1740
           ,x"02e0" -- 1742
           ,x"efa8" -- 1744
           ,x"06a0" -- 1746
           ,x"8094" -- 1748
           ,x"02e0" -- 174A
           ,x"efa8" -- 174C
           ,x"0201" -- 174E
           ,x"c850" -- 1750
           ,x"10e3" -- 1752
           ,x"ef88" -- 1754
           ,x"8158" -- 1756
           ,x"0420" -- 1758
           ,x"8194" -- 175A
           ,x"0380" -- 175C
           ,x"1000" -- 175E
           ,x"0280" -- 1760
           ,x"2000" -- 1762
           ,x"1602" -- 1764
           ,x"0420" -- 1766
           ,x"8198" -- 1768
           ,x"0380" -- 176A
           ,x"eec0" -- 176C
           ,x"81b0" -- 176E
           ,x"eec0" -- 1770
           ,x"81c0" -- 1772
           ,x"eec0" -- 1774
           ,x"81ce" -- 1776
           ,x"eec0" -- 1778
           ,x"81da" -- 177A
           ,x"eec0" -- 177C
           ,x"81d6" -- 177E
           ,x"eec0" -- 1780
           ,x"81e6" -- 1782
           ,x"eec0" -- 1784
           ,x"81e2" -- 1786
           ,x"eec0" -- 1788
           ,x"8228" -- 178A
           ,x"eec0" -- 178C
           ,x"81ac" -- 178E
           ,x"eec0" -- 1790
           ,x"81c8" -- 1792
           ,x"eec0" -- 1794
           ,x"82ac" -- 1796
           ,x"eec0" -- 1798
           ,x"82a8" -- 179A
           ,x"eec0" -- 179C
           ,x"8336" -- 179E
           ,x"eec0" -- 17A0
           ,x"8384" -- 17A2
           ,x"eec0" -- 17A4
           ,x"8330" -- 17A6
           ,x"eec0" -- 17A8
           ,x"837e" -- 17AA
           ,x"c33e" -- 17AC
           ,x"1002" -- 17AE
           ,x"04c4" -- 17B0
           ,x"c31d" -- 17B2
           ,x"020a" -- 17B4
           ,x"edde" -- 17B6
           ,x"024c" -- 17B8
           ,x"ff00" -- 17BA
           ,x"c68c" -- 17BC
           ,x"1015" -- 17BE
           ,x"04c4" -- 17C0
           ,x"020a" -- 17C2
           ,x"c8b9" -- 17C4
           ,x"1011" -- 17C6
           ,x"c32d" -- 17C8
           ,x"000e" -- 17CA
           ,x"771c" -- 17CC
           ,x"04c4" -- 17CE
           ,x"c2a0" -- 17D0
           ,x"ed04" -- 17D2
           ,x"100a" -- 17D4
           ,x"0704" -- 17D6
           ,x"1001" -- 17D8
           ,x"04c4" -- 17DA
           ,x"c2ad" -- 17DC
           ,x"0002" -- 17DE
           ,x"1004" -- 17E0
           ,x"0704" -- 17E2
           ,x"1001" -- 17E4
           ,x"04c4" -- 17E6
           ,x"c2be" -- 17E8
           ,x"06a0" -- 17EA
           ,x"8226" -- 17EC
           ,x"0208" -- 17EE
           ,x"ed40" -- 17F0
           ,x"c1c8" -- 17F2
           ,x"de3a" -- 17F4
           ,x"1309" -- 17F6
           ,x"150f" -- 17F8
           ,x"c104" -- 17FA
           ,x"130d" -- 17FC
           ,x"04cb" -- 17FE
           ,x"0608" -- 1800
           ,x"d2d8" -- 1802
           ,x"050b" -- 1804
           ,x"d60b" -- 1806
           ,x"1001" -- 1808
           ,x"0648" -- 180A
           ,x"81c8" -- 180C
           ,x"1401" -- 180E
           ,x"0588" -- 1810
           ,x"06a0" -- 1812
           ,x"823a" -- 1814
           ,x"0380" -- 1816
           ,x"0288" -- 1818
           ,x"ed8e" -- 181A
           ,x"1aeb" -- 181C
           ,x"0608" -- 181E
           ,x"06a0" -- 1820
           ,x"823a" -- 1822
           ,x"10e2" -- 1824
           ,x"045b" -- 1826
           ,x"c220" -- 1828
           ,x"ed2e" -- 182A
           ,x"0206" -- 182C
           ,x"0600" -- 182E
           ,x"0606" -- 1830
           ,x"16fe" -- 1832
           ,x"0608" -- 1834
           ,x"16fa" -- 1836
           ,x"0380" -- 1838
           ,x"c18b" -- 183A
           ,x"c808" -- 183C
           ,x"eee8" -- 183E
           ,x"c160" -- 1840
           ,x"8044" -- 1842
           ,x"c2e0" -- 1844
           ,x"ed3e" -- 1846
           ,x"1301" -- 1848
           ,x"041b" -- 184A
           ,x"04e0" -- 184C
           ,x"eeee" -- 184E
           ,x"020b" -- 1850
           ,x"8064" -- 1852
           ,x"0202" -- 1854
           ,x"ed90" -- 1856
           ,x"0203" -- 1858
           ,x"0010" -- 185A
           ,x"c33b" -- 185C
           ,x"130e" -- 185E
           ,x"2320" -- 1860
           ,x"b920" -- 1862
           ,x"1611" -- 1864
           ,x"024c" -- 1866
           ,x"7ffe" -- 1868
           ,x"c487" -- 186A
           ,x"0722" -- 186C
           ,x"0002" -- 186E
           ,x"2160" -- 1870
           ,x"b920" -- 1872
           ,x"1603" -- 1874
           ,x"05a0" -- 1876
           ,x"eeee" -- 1878
           ,x"1d13" -- 187A
           ,x"0b15" -- 187C
           ,x"1303" -- 187E
           ,x"8cb2" -- 1880
           ,x"0603" -- 1882
           ,x"16eb" -- 1884
           ,x"0456" -- 1886
           ,x"2160" -- 1888
           ,x"b920" -- 188A
           ,x"16f7" -- 188C
           ,x"c00c" -- 188E
           ,x"c31c" -- 1890
           ,x"cb07" -- 1892
           ,x"0012" -- 1894
           ,x"cb08" -- 1896
           ,x"0014" -- 1898
           ,x"cb02" -- 189A
           ,x"0016" -- 189C
           ,x"0410" -- 189E
           ,x"10ed" -- 18A0
           ,x"6100" -- 18A2
           ,x"7a00" -- 18A4
           ,x"e000" -- 18A6
           ,x"0704" -- 18A8
           ,x"1001" -- 18AA
           ,x"04c4" -- 18AC
           ,x"c80c" -- 18AE
           ,x"8034" -- 18B0
           ,x"020c" -- 18B2
           ,x"0000" -- 18B4
           ,x"1f15" -- 18B6
           ,x"1305" -- 18B8
           ,x"c104" -- 18BA
           ,x"16fc" -- 18BC
           ,x"c320" -- 18BE
           ,x"8034" -- 18C0
           ,x"0380" -- 18C2
           ,x"04dd" -- 18C4
           ,x"361d" -- 18C6
           ,x"1e12" -- 18C8
           ,x"881d" -- 18CA
           ,x"82a2" -- 18CC
           ,x"1a05" -- 18CE
           ,x"881d" -- 18D0
           ,x"82a4" -- 18D2
           ,x"1b02" -- 18D4
           ,x"a760" -- 18D6
           ,x"82a6" -- 18D8
           ,x"c31d" -- 18DA
           ,x"028c" -- 18DC
           ,x"1400" -- 18DE
           ,x"1603" -- 18E0
           ,x"020c" -- 18E2
           ,x"0500" -- 18E4
           ,x"1017" -- 18E6
           ,x"028c" -- 18E8
           ,x"0300" -- 18EA
           ,x"1603" -- 18EC
           ,x"020c" -- 18EE
           ,x"1700" -- 18F0
           ,x"1011" -- 18F2
           ,x"028c" -- 18F4
           ,x"0800" -- 18F6
           ,x"1603" -- 18F8
           ,x"020c" -- 18FA
           ,x"7f00" -- 18FC
           ,x"100b" -- 18FE
           ,x"028c" -- 1900
           ,x"1300" -- 1902
           ,x"1603" -- 1904
           ,x"020c" -- 1906
           ,x"0800" -- 1908
           ,x"1005" -- 190A
           ,x"028c" -- 190C
           ,x"0400" -- 190E
           ,x"1602" -- 1910
           ,x"020c" -- 1912
           ,x"0900" -- 1914
           ,x"c74c" -- 1916
           ,x"c320" -- 1918
           ,x"8034" -- 191A
           ,x"0420" -- 191C
           ,x"8454" -- 191E
           ,x"c104" -- 1920
           ,x"1605" -- 1922
           ,x"981d" -- 1924
           ,x"c84e" -- 1926
           ,x"1601" -- 1928
           ,x"05ce" -- 192A
           ,x"05ce" -- 192C
           ,x"0380" -- 192E
           ,x"c020" -- 1930
           ,x"804c" -- 1932
           ,x"1323" -- 1934
           ,x"d820" -- 1936
           ,x"ed91" -- 1938
           ,x"8348" -- 193A
           ,x"06a0" -- 193C
           ,x"8432" -- 193E
           ,x"0080" -- 1940
           ,x"9081" -- 1942
           ,x"0182" -- 1944
           ,x"0184" -- 1946
           ,x"0087" -- 1948
           ,x"0000" -- 194A
           ,x"0420" -- 194C
           ,x"8bfe" -- 194E
           ,x"0208" -- 1950
           ,x"4400" -- 1952
           ,x"06a0" -- 1954
           ,x"8444" -- 1956
           ,x"020b" -- 1958
           ,x"03c0" -- 195A
           ,x"04e0" -- 195C
           ,x"ef42" -- 195E
           ,x"d820" -- 1960
           ,x"c0e4" -- 1962
           ,x"0000" -- 1964
           ,x"060b" -- 1966
           ,x"16f9" -- 1968
           ,x"d820" -- 196A
           ,x"c0e4" -- 196C
           ,x"ed90" -- 196E
           ,x"04e0" -- 1970
           ,x"804c" -- 1972
           ,x"06a0" -- 1974
           ,x"8432" -- 1976
           ,x"d081" -- 1978
           ,x"0000" -- 197A
           ,x"0380" -- 197C
           ,x"c020" -- 197E
           ,x"804c" -- 1980
           ,x"16fc" -- 1982
           ,x"d820" -- 1984
           ,x"ed91" -- 1986
           ,x"839c" -- 1988
           ,x"06a0" -- 198A
           ,x"8432" -- 198C
           ,x"0280" -- 198E
           ,x"8081" -- 1990
           ,x"0682" -- 1992
           ,x"ff83" -- 1994
           ,x"0384" -- 1996
           ,x"3685" -- 1998
           ,x"0786" -- 199A
           ,x"0087" -- 199C
           ,x"0000" -- 199E
           ,x"04c6" -- 19A0
           ,x"0207" -- 19A2
           ,x"0000" -- 19A4
           ,x"0208" -- 19A6
           ,x"7800" -- 19A8
           ,x"06a0" -- 19AA
           ,x"8444" -- 19AC
           ,x"0208" -- 19AE
           ,x"0800" -- 19B0
           ,x"d5c6" -- 19B2
           ,x"c208" -- 19B4
           ,x"0608" -- 19B6
           ,x"16fc" -- 19B8
           ,x"0208" -- 19BA
           ,x"5b00" -- 19BC
           ,x"06a0" -- 19BE
           ,x"8444" -- 19C0
           ,x"0208" -- 19C2
           ,x"0100" -- 19C4
           ,x"0206" -- 19C6
           ,x"d000" -- 19C8
           ,x"d5c6" -- 19CA
           ,x"c208" -- 19CC
           ,x"0608" -- 19CE
           ,x"16fc" -- 19D0
           ,x"0208" -- 19D2
           ,x"5800" -- 19D4
           ,x"06a0" -- 19D6
           ,x"8444" -- 19D8
           ,x"070b" -- 19DA
           ,x"058b" -- 19DC
           ,x"06cb" -- 19DE
           ,x"d80b" -- 19E0
           ,x"0000" -- 19E2
           ,x"06cb" -- 19E4
           ,x"028b" -- 19E6
           ,x"0300" -- 19E8
           ,x"1af8" -- 19EA
           ,x"0208" -- 19EC
           ,x"4000" -- 19EE
           ,x"06a0" -- 19F0
           ,x"8444" -- 19F2
           ,x"020b" -- 19F4
           ,x"1800" -- 19F6
           ,x"04e0" -- 19F8
           ,x"ef42" -- 19FA
           ,x"d820" -- 19FC
           ,x"c8bb" -- 19FE
           ,x"0000" -- 1A00
           ,x"060b" -- 1A02
           ,x"16f9" -- 1A04
           ,x"0208" -- 1A06
           ,x"6000" -- 1A08
           ,x"06a0" -- 1A0A
           ,x"8444" -- 1A0C
           ,x"020b" -- 1A0E
           ,x"1800" -- 1A10
           ,x"d820" -- 1A12
           ,x"ed91" -- 1A14
           ,x"0000" -- 1A16
           ,x"c208" -- 1A18
           ,x"060b" -- 1A1A
           ,x"16fa" -- 1A1C
           ,x"0720" -- 1A1E
           ,x"804c" -- 1A20
           ,x"d820" -- 1A22
           ,x"8bda" -- 1A24
           ,x"842c" -- 1A26
           ,x"06a0" -- 1A28
           ,x"8432" -- 1A2A
           ,x"c081" -- 1A2C
           ,x"0000" -- 1A2E
           ,x"0380" -- 1A30
           ,x"d83b" -- 1A32
           ,x"0000" -- 1A34
           ,x"86db" -- 1A36
           ,x"d83b" -- 1A38
           ,x"0000" -- 1A3A
           ,x"c6db" -- 1A3C
           ,x"16f9" -- 1A3E
           ,x"05cb" -- 1A40
           ,x"045b" -- 1A42
           ,x"06c8" -- 1A44
           ,x"d808" -- 1A46
           ,x"0000" -- 1A48
           ,x"06c8" -- 1A4A
           ,x"d808" -- 1A4C
           ,x"0000" -- 1A4E
           ,x"86db" -- 1A50
           ,x"045b" -- 1A52
           ,x"eee0" -- 1A54
           ,x"8458" -- 1A56
           ,x"c320" -- 1A58
           ,x"8046" -- 1A5A
           ,x"1610" -- 1A5C
           ,x"c2ed" -- 1A5E
           ,x"001a" -- 1A60
           ,x"981b" -- 1A62
           ,x"c84e" -- 1A64
           ,x"160b" -- 1A66
           ,x"04e0" -- 1A68
           ,x"ed3a" -- 1A6A
           ,x"020e" -- 1A6C
           ,x"8dde" -- 1A6E
           ,x"c320" -- 1A70
           ,x"ede4" -- 1A72
           ,x"1602" -- 1A74
           ,x"020e" -- 1A76
           ,x"8116" -- 1A78
           ,x"020d" -- 1A7A
           ,x"efa8" -- 1A7C
           ,x"0380" -- 1A7E
           ,x"d220" -- 1A80
           ,x"ef43" -- 1A82
           ,x"0988" -- 1A84
           ,x"0228" -- 1A86
           ,x"0007" -- 1A88
           ,x"0938" -- 1A8A
           ,x"d1e0" -- 1A8C
           ,x"ef42" -- 1A8E
           ,x"0987" -- 1A90
           ,x"0227" -- 1A92
           ,x"0007" -- 1A94
           ,x"0937" -- 1A96
           ,x"0287" -- 1A98
           ,x"001f" -- 1A9A
           ,x"1202" -- 1A9C
           ,x"04c7" -- 1A9E
           ,x"0588" -- 1AA0
           ,x"0288" -- 1AA2
           ,x"0017" -- 1AA4
           ,x"1201" -- 1AA6
           ,x"04c8" -- 1AA8
           ,x"0a58" -- 1AAA
           ,x"a207" -- 1AAC
           ,x"0a38" -- 1AAE
           ,x"0228" -- 1AB0
           ,x"4000" -- 1AB2
           ,x"0694" -- 1AB4
           ,x"8289" -- 1AB6
           ,x"1b27" -- 1AB8
           ,x"d039" -- 1ABA
           ,x"9800" -- 1ABC
           ,x"c0e4" -- 1ABE
           ,x"1a34" -- 1AC0
           ,x"0420" -- 1AC2
           ,x"8be0" -- 1AC4
           ,x"0201" -- 1AC6
           ,x"ef48" -- 1AC8
           ,x"0200" -- 1ACA
           ,x"0008" -- 1ACC
           ,x"c080" -- 1ACE
           ,x"a200" -- 1AD0
           ,x"d831" -- 1AD2
           ,x"0000" -- 1AD4
           ,x"0600" -- 1AD6
           ,x"16fc" -- 1AD8
           ,x"0228" -- 1ADA
           ,x"1ff8" -- 1ADC
           ,x"0694" -- 1ADE
           ,x"d820" -- 1AE0
           ,x"ed91" -- 1AE2
           ,x"0000" -- 1AE4
           ,x"0602" -- 1AE6
           ,x"16fb" -- 1AE8
           ,x"0228" -- 1AEA
           ,x"e008" -- 1AEC
           ,x"0694" -- 1AEE
           ,x"0288" -- 1AF0
           ,x"5800" -- 1AF2
           ,x"1ae0" -- 1AF4
           ,x"0228" -- 1AF6
           ,x"e800" -- 1AF8
           ,x"10dc" -- 1AFA
           ,x"04e0" -- 1AFC
           ,x"ed36" -- 1AFE
           ,x"10da" -- 1B00
           ,x"0720" -- 1B02
           ,x"ed36" -- 1B04
           ,x"10d7" -- 1B06
           ,x"0248" -- 1B08
           ,x"1ff8" -- 1B0A
           ,x"06c8" -- 1B0C
           ,x"d808" -- 1B0E
           ,x"ef42" -- 1B10
           ,x"0ab8" -- 1B12
           ,x"d808" -- 1B14
           ,x"ef43" -- 1B16
           ,x"0380" -- 1B18
           ,x"ef00" -- 1B1A
           ,x"851e" -- 1B1C
           ,x"0204" -- 1B1E
           ,x"8444" -- 1B20
           ,x"c020" -- 1B22
           ,x"804c" -- 1B24
           ,x"16ac" -- 1B26
           ,x"102e" -- 1B28
           ,x"06a0" -- 1B2A
           ,x"872c" -- 1B2C
           ,x"0b09" -- 1B2E
           ,x"0f08" -- 1B30
           ,x"180a" -- 1B32
           ,x"1b0b" -- 1B34
           ,x"200c" -- 1B36
           ,x"250d" -- 1B38
           ,x"e71c" -- 1B3A
           ,x"ea1d" -- 1B3C
           ,x"221e" -- 1B3E
           ,x"0000" -- 1B40
           ,x"10b9" -- 1B42
           ,x"0228" -- 1B44
           ,x"0008" -- 1B46
           ,x"0694" -- 1B48
           ,x"10d2" -- 1B4A
           ,x"0228" -- 1B4C
           ,x"fff8" -- 1B4E
           ,x"0694" -- 1B50
           ,x"0288" -- 1B52
           ,x"4000" -- 1B54
           ,x"14af" -- 1B56
           ,x"0228" -- 1B58
           ,x"1800" -- 1B5A
           ,x"10ab" -- 1B5C
           ,x"0228" -- 1B5E
           ,x"0100" -- 1B60
           ,x"10f2" -- 1B62
           ,x"0228" -- 1B64
           ,x"ff00" -- 1B66
           ,x"10f3" -- 1B68
           ,x"c8f2" -- 1B6A
           ,x"83d2" -- 1B6C
           ,x"0420" -- 1B6E
           ,x"856a" -- 1B70
           ,x"0208" -- 1B72
           ,x"4000" -- 1B74
           ,x"109e" -- 1B76
           ,x"0248" -- 1B78
           ,x"ff00" -- 1B7A
           ,x"04e0" -- 1B7C
           ,x"ed34" -- 1B7E
           ,x"1099" -- 1B80
           ,x"c8f2" -- 1B82
           ,x"8336" -- 1B84
           ,x"d1e0" -- 1B86
           ,x"ef43" -- 1B88
           ,x"0987" -- 1B8A
           ,x"39e0" -- 1B8C
           ,x"86e0" -- 1B8E
           ,x"d1e0" -- 1B90
           ,x"ef42" -- 1B92
           ,x"0987" -- 1B94
           ,x"a207" -- 1B96
           ,x"0288" -- 1B98
           ,x"03c0" -- 1B9A
           ,x"1a02" -- 1B9C
           ,x"0420" -- 1B9E
           ,x"8582" -- 1BA0
           ,x"0228" -- 1BA2
           ,x"4400" -- 1BA4
           ,x"c020" -- 1BA6
           ,x"ed36" -- 1BA8
           ,x"1604" -- 1BAA
           ,x"0694" -- 1BAC
           ,x"d820" -- 1BAE
           ,x"ed90" -- 1BB0
           ,x"0000" -- 1BB2
           ,x"0694" -- 1BB4
           ,x"8289" -- 1BB6
           ,x"1b42" -- 1BB8
           ,x"d039" -- 1BBA
           ,x"c820" -- 1BBC
           ,x"8030" -- 1BBE
           ,x"8030" -- 1BC0
           ,x"1603" -- 1BC2
           ,x"9800" -- 1BC4
           ,x"c0e4" -- 1BC6
           ,x"1a76" -- 1BC8
           ,x"d800" -- 1BCA
           ,x"0000" -- 1BCC
           ,x"0588" -- 1BCE
           ,x"0288" -- 1BD0
           ,x"47bf" -- 1BD2
           ,x"12f0" -- 1BD4
           ,x"c820" -- 1BD6
           ,x"8032" -- 1BD8
           ,x"8032" -- 1BDA
           ,x"1303" -- 1BDC
           ,x"0228" -- 1BDE
           ,x"fc40" -- 1BE0
           ,x"10e8" -- 1BE2
           ,x"c1c8" -- 1BE4
           ,x"0227" -- 1BE6
           ,x"ffd8" -- 1BE8
           ,x"0208" -- 1BEA
           ,x"0428" -- 1BEC
           ,x"0694" -- 1BEE
           ,x"04c1" -- 1BF0
           ,x"d860" -- 1BF2
           ,x"0000" -- 1BF4
           ,x"c8f2" -- 1BF6
           ,x"0581" -- 1BF8
           ,x"0281" -- 1BFA
           ,x"0398" -- 1BFC
           ,x"1af9" -- 1BFE
           ,x"0208" -- 1C00
           ,x"4400" -- 1C02
           ,x"0694" -- 1C04
           ,x"04c1" -- 1C06
           ,x"d821" -- 1C08
           ,x"c8f2" -- 1C0A
           ,x"0000" -- 1C0C
           ,x"0581" -- 1C0E
           ,x"0281" -- 1C10
           ,x"0398" -- 1C12
           ,x"1af9" -- 1C14
           ,x"0201" -- 1C16
           ,x"0028" -- 1C18
           ,x"d820" -- 1C1A
           ,x"c0e4" -- 1C1C
           ,x"0000" -- 1C1E
           ,x"d820" -- 1C20
           ,x"c0e4" -- 1C22
           ,x"0000" -- 1C24
           ,x"0641" -- 1C26
           ,x"16f8" -- 1C28
           ,x"c207" -- 1C2A
           ,x"0694" -- 1C2C
           ,x"10c3" -- 1C2E
           ,x"0288" -- 1C30
           ,x"4400" -- 1C32
           ,x"14c0" -- 1C34
           ,x"0228" -- 1C36
           ,x"03c0" -- 1C38
           ,x"0694" -- 1C3A
           ,x"10bc" -- 1C3C
           ,x"0228" -- 1C3E
           ,x"c000" -- 1C40
           ,x"0694" -- 1C42
           ,x"04c3" -- 1C44
           ,x"d0e0" -- 1C46
           ,x"0000" -- 1C48
           ,x"0228" -- 1C4A
           ,x"4000" -- 1C4C
           ,x"0694" -- 1C4E
           ,x"c060" -- 1C50
           ,x"ed36" -- 1C52
           ,x"1603" -- 1C54
           ,x"d820" -- 1C56
           ,x"c84b" -- 1C58
           ,x"0000" -- 1C5A
           ,x"0228" -- 1C5C
           ,x"bc00" -- 1C5E
           ,x"04c7" -- 1C60
           ,x"3de0" -- 1C62
           ,x"86e0" -- 1C64
           ,x"02a1" -- 1C66
           ,x"d821" -- 1C68
           ,x"000f" -- 1C6A
           ,x"ef43" -- 1C6C
           ,x"d821" -- 1C6E
           ,x"0011" -- 1C70
           ,x"ef42" -- 1C72
           ,x"d803" -- 1C74
           ,x"ed90" -- 1C76
           ,x"0953" -- 1C78
           ,x"c203" -- 1C7A
           ,x"0228" -- 1C7C
           ,x"0800" -- 1C7E
           ,x"0694" -- 1C80
           ,x"0208" -- 1C82
           ,x"ef48" -- 1C84
           ,x"c048" -- 1C86
           ,x"0207" -- 1C88
           ,x"0008" -- 1C8A
           ,x"c087" -- 1C8C
           ,x"de20" -- 1C8E
           ,x"0000" -- 1C90
           ,x"0607" -- 1C92
           ,x"16fc" -- 1C94
           ,x"0208" -- 1C96
           ,x"4bf8" -- 1C98
           ,x"0694" -- 1C9A
           ,x"d031" -- 1C9C
           ,x"0540" -- 1C9E
           ,x"d800" -- 1CA0
           ,x"0000" -- 1CA2
           ,x"0602" -- 1CA4
           ,x"16fa" -- 1CA6
           ,x"0380" -- 1CA8
           ,x"04e0" -- 1CAA
           ,x"ed36" -- 1CAC
           ,x"10c6" -- 1CAE
           ,x"0720" -- 1CB0
           ,x"ed36" -- 1CB2
           ,x"10c3" -- 1CB4
           ,x"06a0" -- 1CB6
           ,x"872c" -- 1CB8
           ,x"0b09" -- 1CBA
           ,x"0f08" -- 1CBC
           ,x"120a" -- 1CBE
           ,x"150b" -- 1CC0
           ,x"180c" -- 1CC2
           ,x"260d" -- 1CC4
           ,x"f81c" -- 1CC6
           ,x"fb1d" -- 1CC8
           ,x"221e" -- 1CCA
           ,x"0000" -- 1CCC
           ,x"10b6" -- 1CCE
           ,x"0588" -- 1CD0
           ,x"0694" -- 1CD2
           ,x"0460" -- 1CD4
           ,x"85d0" -- 1CD6
           ,x"0608" -- 1CD8
           ,x"0694" -- 1CDA
           ,x"10a9" -- 1CDC
           ,x"0228" -- 1CDE
           ,x"0028" -- 1CE0
           ,x"10f7" -- 1CE2
           ,x"0228" -- 1CE4
           ,x"ffd8" -- 1CE6
           ,x"10f8" -- 1CE8
           ,x"0208" -- 1CEA
           ,x"4400" -- 1CEC
           ,x"0694" -- 1CEE
           ,x"0201" -- 1CF0
           ,x"03c0" -- 1CF2
           ,x"c820" -- 1CF4
           ,x"c0e4" -- 1CF6
           ,x"0000" -- 1CF8
           ,x"0601" -- 1CFA
           ,x"16fb" -- 1CFC
           ,x"0208" -- 1CFE
           ,x"4400" -- 1D00
           ,x"0694" -- 1D02
           ,x"10e4" -- 1D04
           ,x"0228" -- 1D06
           ,x"bc00" -- 1D08
           ,x"04c7" -- 1D0A
           ,x"3de0" -- 1D0C
           ,x"86e0" -- 1D0E
           ,x"39e0" -- 1D10
           ,x"86e0" -- 1D12
           ,x"0228" -- 1D14
           ,x"4400" -- 1D16
           ,x"04e0" -- 1D18
           ,x"ed34" -- 1D1A
           ,x"10f2" -- 1D1C
           ,x"0420" -- 1D1E
           ,x"8d70" -- 1D20
           ,x"0032" -- 1D22
           ,x"04c0" -- 1D24
           ,x"d038" -- 1D26
           ,x"c800" -- 1D28
           ,x"ede8" -- 1D2A
           ,x"c08b" -- 1D2C
           ,x"04c1" -- 1D2E
           ,x"d07b" -- 1D30
           ,x"1305" -- 1D32
           ,x"9ec0" -- 1D34
           ,x"16fc" -- 1D36
           ,x"0871" -- 1D38
           ,x"a081" -- 1D3A
           ,x"0452" -- 1D3C
           ,x"058b" -- 1D3E
           ,x"045b" -- 1D40
           ,x"0420" -- 1D42
           ,x"8d70" -- 1D44
           ,x"0032" -- 1D46
           ,x"0420" -- 1D48
           ,x"8d70" -- 1D4A
           ,x"0032" -- 1D4C
           ,x"0420" -- 1D4E
           ,x"8d70" -- 1D50
           ,x"0032" -- 1D52
           ,x"0420" -- 1D54
           ,x"8194" -- 1D56
           ,x"10fd" -- 1D58
           ,x"1001" -- 1D5A
           ,x"100b" -- 1D5C
           ,x"0420" -- 1D5E
           ,x"816c" -- 1D60
           ,x"0280" -- 1D62
           ,x"5900" -- 1D64
           ,x"1304" -- 1D66
           ,x"0280" -- 1D68
           ,x"4e00" -- 1D6A
           ,x"1602" -- 1D6C
           ,x"05cb" -- 1D6E
           ,x"05cb" -- 1D70
           ,x"045b" -- 1D72
           ,x"0460" -- 1D74
           ,x"8116" -- 1D76
           ,x"06a0" -- 1D78
           ,x"c4d0" -- 1D7A
           ,x"1077" -- 1D7C
           ,x"04c1" -- 1D7E
           ,x"d052" -- 1D80
           ,x"04c4" -- 1D82
           ,x"c0a0" -- 1D84
           ,x"ef68" -- 1D86
           ,x"60a0" -- 1D88
           ,x"887e" -- 1D8A
           ,x"1110" -- 1D8C
           ,x"c820" -- 1D8E
           ,x"8012" -- 1D90
           ,x"ef7e" -- 1D92
           ,x"0420" -- 1D94
           ,x"bc32" -- 1D96
           ,x"c820" -- 1D98
           ,x"88ca" -- 1D9A
           ,x"ef7e" -- 1D9C
           ,x"0420" -- 1D9E
           ,x"bc3e" -- 1DA0
           ,x"c820" -- 1DA2
           ,x"8012" -- 1DA4
           ,x"ef7e" -- 1DA6
           ,x"0420" -- 1DA8
           ,x"beac" -- 1DAA
           ,x"0584" -- 1DAC
           ,x"c820" -- 1DAE
           ,x"8012" -- 1DB0
           ,x"ef7e" -- 1DB2
           ,x"0420" -- 1DB4
           ,x"bc32" -- 1DB6
           ,x"c820" -- 1DB8
           ,x"88c2" -- 1DBA
           ,x"ef7e" -- 1DBC
           ,x"0420" -- 1DBE
           ,x"bc4e" -- 1DC0
           ,x"c0a0" -- 1DC2
           ,x"ef68" -- 1DC4
           ,x"c820" -- 1DC6
           ,x"8012" -- 1DC8
           ,x"ef7e" -- 1DCA
           ,x"0420" -- 1DCC
           ,x"bc3e" -- 1DCE
           ,x"c082" -- 1DD0
           ,x"111e" -- 1DD2
           ,x"c820" -- 1DD4
           ,x"88c4" -- 1DD6
           ,x"ef7e" -- 1DD8
           ,x"0420" -- 1DDA
           ,x"bc4a" -- 1DDC
           ,x"c820" -- 1DDE
           ,x"8000" -- 1DE0
           ,x"ef7e" -- 1DE2
           ,x"0420" -- 1DE4
           ,x"bc32" -- 1DE6
           ,x"c820" -- 1DE8
           ,x"8012" -- 1DEA
           ,x"ef7e" -- 1DEC
           ,x"0420" -- 1DEE
           ,x"bc3e" -- 1DF0
           ,x"c820" -- 1DF2
           ,x"88c4" -- 1DF4
           ,x"ef7e" -- 1DF6
           ,x"0420" -- 1DF8
           ,x"bd84" -- 1DFA
           ,x"c820" -- 1DFC
           ,x"88ca" -- 1DFE
           ,x"ef7e" -- 1E00
           ,x"0420" -- 1E02
           ,x"bc4e" -- 1E04
           ,x"c820" -- 1E06
           ,x"8000" -- 1E08
           ,x"ef7e" -- 1E0A
           ,x"0420" -- 1E0C
           ,x"beac" -- 1E0E
           ,x"c820" -- 1E10
           ,x"8000" -- 1E12
           ,x"ef7e" -- 1E14
           ,x"0420" -- 1E16
           ,x"bc32" -- 1E18
           ,x"06a0" -- 1E1A
           ,x"c4f4" -- 1E1C
           ,x"887c" -- 1E1E
           ,x"c820" -- 1E20
           ,x"8002" -- 1E22
           ,x"ef7e" -- 1E24
           ,x"0420" -- 1E26
           ,x"bc32" -- 1E28
           ,x"06a0" -- 1E2A
           ,x"c512" -- 1E2C
           ,x"889c" -- 1E2E
           ,x"c820" -- 1E30
           ,x"8002" -- 1E32
           ,x"ef7e" -- 1E34
           ,x"0420" -- 1E36
           ,x"beac" -- 1E38
           ,x"c820" -- 1E3A
           ,x"8000" -- 1E3C
           ,x"ef7e" -- 1E3E
           ,x"0420" -- 1E40
           ,x"bd84" -- 1E42
           ,x"c082" -- 1E44
           ,x"1105" -- 1E46
           ,x"c820" -- 1E48
           ,x"88c6" -- 1E4A
           ,x"ef7e" -- 1E4C
           ,x"0420" -- 1E4E
           ,x"bc4a" -- 1E50
           ,x"0604" -- 1E52
           ,x"1605" -- 1E54
           ,x"c820" -- 1E56
           ,x"88c8" -- 1E58
           ,x"ef7e" -- 1E5A
           ,x"0420" -- 1E5C
           ,x"bc4a" -- 1E5E
           ,x"0b13" -- 1E60
           ,x"4820" -- 1E62
           ,x"bfca" -- 1E64
           ,x"ef68" -- 1E66
           ,x"a803" -- 1E68
           ,x"ef68" -- 1E6A
           ,x"0460" -- 1E6C
           ,x"b6be" -- 1E6E
           ,x"4044" -- 1E70
           ,x"9851" -- 1E72
           ,x"7a7b" -- 1E74
           ,x"411b" -- 1E76
           ,x"b67a" -- 1E78
           ,x"e858" -- 1E7A
           ,x"0004" -- 1E7C
           ,x"4110" -- 1E7E
           ,x"0000" -- 1E80
           ,x"0000" -- 1E82
           ,x"4225" -- 1E84
           ,x"10eb" -- 1E86
           ,x"4200" -- 1E88
           ,x"42cf" -- 1E8A
           ,x"b153" -- 1E8C
           ,x"9710" -- 1E8E
           ,x"4316" -- 1E90
           ,x"ca99" -- 1E92
           ,x"3433" -- 1E94
           ,x"42c5" -- 1E96
           ,x"33fe" -- 1E98
           ,x"142d" -- 1E9A
           ,x"0003" -- 1E9C
           ,x"41c9" -- 1E9E
           ,x"8867" -- 1EA0
           ,x"f42a" -- 1EA2
           ,x"427d" -- 1EA4
           ,x"9444" -- 1EA6
           ,x"406e" -- 1EA8
           ,x"4312" -- 1EAA
           ,x"aed9" -- 1EAC
           ,x"3e72" -- 1EAE
           ,x"42c5" -- 1EB0
           ,x"33fe" -- 1EB2
           ,x"142d" -- 1EB4
           ,x"4086" -- 1EB6
           ,x"0a91" -- 1EB8
           ,x"c16c" -- 1EBA
           ,x"c119" -- 1EBC
           ,x"21fb" -- 1EBE
           ,x"5444" -- 1EC0
           ,x"8870" -- 1EC2
           ,x"8876" -- 1EC4
           ,x"88b6" -- 1EC6
           ,x"88bc" -- 1EC8
           ,x"887e" -- 1ECA
           ,x"c820" -- 1ECC
           ,x"801a" -- 1ECE
           ,x"ef9e" -- 1ED0
           ,x"0420" -- 1ED2
           ,x"b558" -- 1ED4
           ,x"c020" -- 1ED6
           ,x"804c" -- 1ED8
           ,x"1612" -- 1EDA
           ,x"0281" -- 1EDC
           ,x"03c0" -- 1EDE
           ,x"1478" -- 1EE0
           ,x"0420" -- 1EE2
           ,x"b526" -- 1EE4
           ,x"c3c8" -- 1EE6
           ,x"c201" -- 1EE8
           ,x"0228" -- 1EEA
           ,x"0400" -- 1EEC
           ,x"06a0" -- 1EEE
           ,x"8444" -- 1EF0
           ,x"04f2" -- 1EF2
           ,x"04f2" -- 1EF4
           ,x"04d2" -- 1EF6
           ,x"d8a0" -- 1EF8
           ,x"0000" -- 1EFA
           ,x"ffff" -- 1EFC
           ,x"1067" -- 1EFE
           ,x"0281" -- 1F00
           ,x"0300" -- 1F02
           ,x"1466" -- 1F04
           ,x"c820" -- 1F06
           ,x"801c" -- 1F08
           ,x"ef9e" -- 1F0A
           ,x"0420" -- 1F0C
           ,x"b558" -- 1F0E
           ,x"c3c8" -- 1F10
           ,x"c201" -- 1F12
           ,x"0a38" -- 1F14
           ,x"06a0" -- 1F16
           ,x"8444" -- 1F18
           ,x"0203" -- 1F1A
           ,x"ef48" -- 1F1C
           ,x"c103" -- 1F1E
           ,x"0200" -- 1F20
           ,x"0008" -- 1F22
           ,x"dce0" -- 1F24
           ,x"0000" -- 1F26
           ,x"0600" -- 1F28
           ,x"16fc" -- 1F2A
           ,x"c202" -- 1F2C
           ,x"0a38" -- 1F2E
           ,x"0228" -- 1F30
           ,x"7800" -- 1F32
           ,x"06a0" -- 1F34
           ,x"8444" -- 1F36
           ,x"0200" -- 1F38
           ,x"0008" -- 1F3A
           ,x"d834" -- 1F3C
           ,x"0000" -- 1F3E
           ,x"0600" -- 1F40
           ,x"16fc" -- 1F42
           ,x"1044" -- 1F44
           ,x"c820" -- 1F46
           ,x"801a" -- 1F48
           ,x"ef9e" -- 1F4A
           ,x"0420" -- 1F4C
           ,x"b558" -- 1F4E
           ,x"c820" -- 1F50
           ,x"801c" -- 1F52
           ,x"ef9e" -- 1F54
           ,x"0420" -- 1F56
           ,x"b558" -- 1F58
           ,x"d082" -- 1F5A
           ,x"163a" -- 1F5C
           ,x"c3c8" -- 1F5E
           ,x"c020" -- 1F60
           ,x"804c" -- 1F62
           ,x"160c" -- 1F64
           ,x"0281" -- 1F66
           ,x"03c0" -- 1F68
           ,x"1433" -- 1F6A
           ,x"c201" -- 1F6C
           ,x"0228" -- 1F6E
           ,x"4400" -- 1F70
           ,x"06a0" -- 1F72
           ,x"8444" -- 1F74
           ,x"06c2" -- 1F76
           ,x"d802" -- 1F78
           ,x"0000" -- 1F7A
           ,x"1028" -- 1F7C
           ,x"0281" -- 1F7E
           ,x"0300" -- 1F80
           ,x"1427" -- 1F82
           ,x"c202" -- 1F84
           ,x"0a38" -- 1F86
           ,x"0228" -- 1F88
           ,x"3800" -- 1F8A
           ,x"06a0" -- 1F8C
           ,x"8444" -- 1F8E
           ,x"0208" -- 1F90
           ,x"0008" -- 1F92
           ,x"c0c8" -- 1F94
           ,x"0200" -- 1F96
           ,x"ef48" -- 1F98
           ,x"c100" -- 1F9A
           ,x"dc20" -- 1F9C
           ,x"0000" -- 1F9E
           ,x"0608" -- 1FA0
           ,x"16fc" -- 1FA2
           ,x"c201" -- 1FA4
           ,x"0a38" -- 1FA6
           ,x"0228" -- 1FA8
           ,x"4000" -- 1FAA
           ,x"06a0" -- 1FAC
           ,x"8444" -- 1FAE
           ,x"d834" -- 1FB0
           ,x"0000" -- 1FB2
           ,x"0603" -- 1FB4
           ,x"16fc" -- 1FB6
           ,x"0228" -- 1FB8
           ,x"2000" -- 1FBA
           ,x"06a0" -- 1FBC
           ,x"8444" -- 1FBE
           ,x"0205" -- 1FC0
           ,x"0008" -- 1FC2
           ,x"d820" -- 1FC4
           ,x"ed91" -- 1FC6
           ,x"0000" -- 1FC8
           ,x"0605" -- 1FCA
           ,x"16fb" -- 1FCC
           ,x"c20f" -- 1FCE
           ,x"1028" -- 1FD0
           ,x"1073" -- 1FD2
           ,x"0420" -- 1FD4
           ,x"819c" -- 1FD6
           ,x"0460" -- 1FD8
           ,x"aef8" -- 1FDA
           ,x"0420" -- 1FDC
           ,x"81a0" -- 1FDE
           ,x"10fb" -- 1FE0
           ,x"06a0" -- 1FE2
           ,x"b52a" -- 1FE4
           ,x"101f" -- 1FE6
           ,x"c820" -- 1FE8
           ,x"8022" -- 1FEA
           ,x"ef9e" -- 1FEC
           ,x"0420" -- 1FEE
           ,x"b558" -- 1FF0
           ,x"0285" -- 1FF2
           ,x"00ff" -- 1FF4
           ,x"1b63" -- 1FF6
           ,x"0204" -- 1FF8
           ,x"0003" -- 1FFA
           ,x"02a6" -- 1FFC
           ,x"05c6" -- 1FFE
           ,x"0280" -- 2000
           ,x"3f00" -- 2002
           ,x"165e" -- 2004
           ,x"c806" -- 2006
           ,x"ef9e" -- 2008
           ,x"05c6" -- 200A
           ,x"0420" -- 200C
           ,x"b558" -- 200E
           ,x"0604" -- 2010
           ,x"16f6" -- 2012
           ,x"3960" -- 2014
           ,x"8c40" -- 2016
           ,x"0226" -- 2018
           ,x"d0ba" -- 201A
           ,x"cd81" -- 201C
           ,x"cd82" -- 201E
           ,x"cd83" -- 2020
           ,x"0608" -- 2022
           ,x"10d9" -- 2024
           ,x"0201" -- 2026
           ,x"d6ba" -- 2028
           ,x"0202" -- 202A
           ,x"d0ba" -- 202C
           ,x"ccb1" -- 202E
           ,x"0282" -- 2030
           ,x"d4b0" -- 2032
           ,x"1afc" -- 2034
           ,x"10d0" -- 2036
           ,x"06a0" -- 2038
           ,x"b52a" -- 203A
           ,x"101f" -- 203C
           ,x"d060" -- 203E
           ,x"ed91" -- 2040
           ,x"06c1" -- 2042
           ,x"c820" -- 2044
           ,x"801c" -- 2046
           ,x"ef9e" -- 2048
           ,x"0420" -- 204A
           ,x"b558" -- 204C
           ,x"0280" -- 204E
           ,x"3f00" -- 2050
           ,x"1605" -- 2052
           ,x"c820" -- 2054
           ,x"801a" -- 2056
           ,x"ef9e" -- 2058
           ,x"0420" -- 205A
           ,x"b558" -- 205C
           ,x"0b41" -- 205E
           ,x"d081" -- 2060
           ,x"0b42" -- 2062
           ,x"d802" -- 2064
           ,x"ed91" -- 2066
           ,x"c060" -- 2068
           ,x"804c" -- 206A
           ,x"16da" -- 206C
           ,x"d802" -- 206E
           ,x"8a76" -- 2070
           ,x"06a0" -- 2072
           ,x"8432" -- 2074
           ,x"0087" -- 2076
           ,x"0000" -- 2078
           ,x"10d3" -- 207A
           ,x"0202" -- 207C
           ,x"1300" -- 207E
           ,x"0588" -- 2080
           ,x"10f0" -- 2082
           ,x"0420" -- 2084
           ,x"81a8" -- 2086
           ,x"c0e0" -- 2088
           ,x"ef42" -- 208A
           ,x"c281" -- 208C
           ,x"06a0" -- 208E
           ,x"bbd6" -- 2090
           ,x"028a" -- 2092
           ,x"00c0" -- 2094
           ,x"140e" -- 2096
           ,x"0281" -- 2098
           ,x"0100" -- 209A
           ,x"140b" -- 209C
           ,x"06c1" -- 209E
           ,x"d281" -- 20A0
           ,x"c80a" -- 20A2
           ,x"ef42" -- 20A4
           ,x"0420" -- 20A6
           ,x"8c5e" -- 20A8
           ,x"ef6b" -- 20AA
           ,x"c803" -- 20AC
           ,x"ef42" -- 20AE
           ,x"0460" -- 20B0
           ,x"b6be" -- 20B2
           ,x"0720" -- 20B4
           ,x"ef6a" -- 20B6
           ,x"10fb" -- 20B8
           ,x"0460" -- 20BA
           ,x"9b68" -- 20BC
           ,x"0460" -- 20BE
           ,x"93fc" -- 20C0
           ,x"0460" -- 20C2
           ,x"aef2" -- 20C4
           ,x"06a0" -- 20C6
           ,x"b52a" -- 20C8
           ,x"1008" -- 20CA
           ,x"c820" -- 20CC
           ,x"8004" -- 20CE
           ,x"ef9e" -- 20D0
           ,x"0420" -- 20D2
           ,x"b558" -- 20D4
           ,x"0420" -- 20D6
           ,x"8188" -- 20D8
           ,x"10a3" -- 20DA
           ,x"0460" -- 20DC
           ,x"89d8" -- 20DE
           ,x"0420" -- 20E0
           ,x"81a8" -- 20E2
           ,x"c820" -- 20E4
           ,x"801a" -- 20E6
           ,x"ef9e" -- 20E8
           ,x"0420" -- 20EA
           ,x"b558" -- 20EC
           ,x"d041" -- 20EE
           ,x"16e4" -- 20F0
           ,x"0a31" -- 20F2
           ,x"0221" -- 20F4
           ,x"7800" -- 20F6
           ,x"c088" -- 20F8
           ,x"c201" -- 20FA
           ,x"06a0" -- 20FC
           ,x"8444" -- 20FE
           ,x"c202" -- 2100
           ,x"0203" -- 2102
           ,x"0004" -- 2104
           ,x"0280" -- 2106
           ,x"3f00" -- 2108
           ,x"16db" -- 210A
           ,x"c820" -- 210C
           ,x"801a" -- 210E
           ,x"ef9e" -- 2110
           ,x"0420" -- 2112
           ,x"b558" -- 2114
           ,x"d801" -- 2116
           ,x"0000" -- 2118
           ,x"06c1" -- 211A
           ,x"d801" -- 211C
           ,x"0000" -- 211E
           ,x"0603" -- 2120
           ,x"16f1" -- 2122
           ,x"0460" -- 2124
           ,x"8a22" -- 2126
           ,x"0420" -- 2128
           ,x"81a8" -- 212A
           ,x"c820" -- 212C
           ,x"802a" -- 212E
           ,x"ef9e" -- 2130
           ,x"0420" -- 2132
           ,x"b558" -- 2134
           ,x"c388" -- 2136
           ,x"028f" -- 2138
           ,x"001f" -- 213A
           ,x"1bbe" -- 213C
           ,x"0a2f" -- 213E
           ,x"022f" -- 2140
           ,x"1b02" -- 2142
           ,x"c20f" -- 2144
           ,x"06a0" -- 2146
           ,x"8444" -- 2148
           ,x"d0a0" -- 214A
           ,x"0000" -- 214C
           ,x"06c2" -- 214E
           ,x"0228" -- 2150
           ,x"3ffe" -- 2152
           ,x"d0a0" -- 2154
           ,x"0000" -- 2156
           ,x"06a0" -- 2158
           ,x"8444" -- 215A
           ,x"c20e" -- 215C
           ,x"c820" -- 215E
           ,x"801a" -- 2160
           ,x"ef9e" -- 2162
           ,x"0420" -- 2164
           ,x"b558" -- 2166
           ,x"c820" -- 2168
           ,x"801e" -- 216A
           ,x"ef9e" -- 216C
           ,x"0420" -- 216E
           ,x"b558" -- 2170
           ,x"06c3" -- 2172
           ,x"d043" -- 2174
           ,x"0280" -- 2176
           ,x"3f00" -- 2178
           ,x"160c" -- 217A
           ,x"c820" -- 217C
           ,x"801c" -- 217E
           ,x"ef9e" -- 2180
           ,x"0420" -- 2182
           ,x"b558" -- 2184
           ,x"c820" -- 2186
           ,x"801e" -- 2188
           ,x"ef9e" -- 218A
           ,x"0420" -- 218C
           ,x"b558" -- 218E
           ,x"06c3" -- 2190
           ,x"d083" -- 2192
           ,x"06c2" -- 2194
           ,x"02a3" -- 2196
           ,x"05c3" -- 2198
           ,x"0204" -- 219A
           ,x"0004" -- 219C
           ,x"d833" -- 219E
           ,x"0000" -- 21A0
           ,x"0604" -- 21A2
           ,x"16fc" -- 21A4
           ,x"10be" -- 21A6
           ,x"0420" -- 21A8
           ,x"81a8" -- 21AA
           ,x"c820" -- 21AC
           ,x"801c" -- 21AE
           ,x"ef9e" -- 21B0
           ,x"0420" -- 21B2
           ,x"b558" -- 21B4
           ,x"c820" -- 21B6
           ,x"801a" -- 21B8
           ,x"ef9e" -- 21BA
           ,x"0420" -- 21BC
           ,x"b558" -- 21BE
           ,x"0203" -- 21C0
           ,x"00c0" -- 21C2
           ,x"c041" -- 21C4
           ,x"1301" -- 21C6
           ,x"05c3" -- 21C8
           ,x"c082" -- 21CA
           ,x"1301" -- 21CC
           ,x"0583" -- 21CE
           ,x"06c3" -- 21D0
           ,x"d803" -- 21D2
           ,x"8bda" -- 21D4
           ,x"06a0" -- 21D6
           ,x"8432" -- 21D8
           ,x"c081" -- 21DA
           ,x"0000" -- 21DC
           ,x"10a2" -- 21DE
           ,x"ef20" -- 21E0
           ,x"8be4" -- 21E2
           ,x"0208" -- 21E4
           ,x"ef48" -- 21E6
           ,x"0209" -- 21E8
           ,x"0001" -- 21EA
           ,x"c2dd" -- 21EC
           ,x"098b" -- 21EE
           ,x"3ae0" -- 21F0
           ,x"8c40" -- 21F2
           ,x"022c" -- 21F4
           ,x"d0ba" -- 21F6
           ,x"020a" -- 21F8
           ,x"0008" -- 21FA
           ,x"101a" -- 21FC
           ,x"ef20" -- 21FE
           ,x"8c02" -- 2200
           ,x"0208" -- 2202
           ,x"4400" -- 2204
           ,x"06a0" -- 2206
           ,x"8444" -- 2208
           ,x"0709" -- 220A
           ,x"0589" -- 220C
           ,x"06c9" -- 220E
           ,x"d809" -- 2210
           ,x"0000" -- 2212
           ,x"06c9" -- 2214
           ,x"0289" -- 2216
           ,x"03c0" -- 2218
           ,x"1af8" -- 221A
           ,x"0208" -- 221C
           ,x"4800" -- 221E
           ,x"06a0" -- 2220
           ,x"8444" -- 2222
           ,x"0208" -- 2224
           ,x"0000" -- 2226
           ,x"04c9" -- 2228
           ,x"020c" -- 222A
           ,x"d0ba" -- 222C
           ,x"020a" -- 222E
           ,x"0800" -- 2230
           ,x"0207" -- 2232
           ,x"0101" -- 2234
           ,x"0706" -- 2236
           ,x"04c5" -- 2238
           ,x"0204" -- 223A
           ,x"0001" -- 223C
           ,x"0203" -- 223E
           ,x"0006" -- 2240
           ,x"0b14" -- 2242
           ,x"0b17" -- 2244
           ,x"1701" -- 2246
           ,x"d1bc" -- 2248
           ,x"2187" -- 224A
           ,x"1601" -- 224C
           ,x"b144" -- 224E
           ,x"0603" -- 2250
           ,x"15f7" -- 2252
           ,x"d605" -- 2254
           ,x"a209" -- 2256
           ,x"060a" -- 2258
           ,x"15ee" -- 225A
           ,x"0380" -- 225C
           ,x"ef40" -- 225E
           ,x"8c62" -- 2260
           ,x"020c" -- 2262
           ,x"2009" -- 2264
           ,x"1009" -- 2266
           ,x"ef40" -- 2268
           ,x"8c6c" -- 226A
           ,x"020c" -- 226C
           ,x"5009" -- 226E
           ,x"1004" -- 2270
           ,x"ef40" -- 2272
           ,x"8c76" -- 2274
           ,x"020c" -- 2276
           ,x"f009" -- 2278
           ,x"d241" -- 227A
           ,x"0989" -- 227C
           ,x"c201" -- 227E
           ,x"0a28" -- 2280
           ,x"0248" -- 2282
           ,x"03e0" -- 2284
           ,x"0288" -- 2286
           ,x"0300" -- 2288
           ,x"142c" -- 228A
           ,x"c281" -- 228C
           ,x"024a" -- 228E
           ,x"0007" -- 2290
           ,x"c009" -- 2292
           ,x"0240" -- 2294
           ,x"0007" -- 2296
           ,x"0939" -- 2298
           ,x"a209" -- 229A
           ,x"0a38" -- 229C
           ,x"a20a" -- 229E
           ,x"06a0" -- 22A0
           ,x"8444" -- 22A2
           ,x"04c9" -- 22A4
           ,x"0220" -- 22A6
           ,x"8d02" -- 22A8
           ,x"d250" -- 22AA
           ,x"d020" -- 22AC
           ,x"0000" -- 22AE
           ,x"0268" -- 22B0
           ,x"4000" -- 22B2
           ,x"06a0" -- 22B4
           ,x"8444" -- 22B6
           ,x"048c" -- 22B8
           ,x"02c9" -- 22BA
           ,x"880c" -- 22BC
           ,x"8c64" -- 22BE
           ,x"1612" -- 22C0
           ,x"0248" -- 22C2
           ,x"bfff" -- 22C4
           ,x"0228" -- 22C6
           ,x"2000" -- 22C8
           ,x"06a0" -- 22CA
           ,x"8444" -- 22CC
           ,x"8f3c" -- 22CE
           ,x"d220" -- 22D0
           ,x"ed91" -- 22D2
           ,x"2260" -- 22D4
           ,x"c0e4" -- 22D6
           ,x"1601" -- 22D8
           ,x"0948" -- 22DA
           ,x"0248" -- 22DC
           ,x"0f00" -- 22DE
           ,x"c27e" -- 22E0
           ,x"d648" -- 22E2
           ,x"0380" -- 22E4
           ,x"d800" -- 22E6
           ,x"0000" -- 22E8
           ,x"880c" -- 22EA
           ,x"8c6e" -- 22EC
           ,x"13fa" -- 22EE
           ,x"0228" -- 22F0
           ,x"2000" -- 22F2
           ,x"06a0" -- 22F4
           ,x"8444" -- 22F6
           ,x"8f3c" -- 22F8
           ,x"d820" -- 22FA
           ,x"ed91" -- 22FC
           ,x"0000" -- 22FE
           ,x"0380" -- 2300
           ,x"8040" -- 2302
           ,x"2010" -- 2304
           ,x"0804" -- 2306
           ,x"0201" -- 2308
           ,x"c80b" -- 230A
           ,x"ed2c" -- 230C
           ,x"0420" -- 230E
           ,x"8184" -- 2310
           ,x"c8d4" -- 2312
           ,x"04e0" -- 2314
           ,x"8046" -- 2316
           ,x"c003" -- 2318
           ,x"06c0" -- 231A
           ,x"0240" -- 231C
           ,x"000f" -- 231E
           ,x"3820" -- 2320
           ,x"9a88" -- 2322
           ,x"c283" -- 2324
           ,x"024a" -- 2326
           ,x"000f" -- 2328
           ,x"a04a" -- 232A
           ,x"c2a0" -- 232C
           ,x"ede4" -- 232E
           ,x"1305" -- 2330
           ,x"c081" -- 2332
           ,x"0420" -- 2334
           ,x"818c" -- 2336
           ,x"0d00" -- 2338
           ,x"101d" -- 233A
           ,x"0281" -- 233C
           ,x"0033" -- 233E
           ,x"1203" -- 2340
           ,x"0202" -- 2342
           ,x"cce0" -- 2344
           ,x"1003" -- 2346
           ,x"a041" -- 2348
           ,x"c0a1" -- 234A
           ,x"8e54" -- 234C
           ,x"0207" -- 234E
           ,x"ee0c" -- 2350
           ,x"06a0" -- 2352
           ,x"8e20" -- 2354
           ,x"75d7" -- 2356
           ,x"0420" -- 2358
           ,x"8180" -- 235A
           ,x"ee0c" -- 235C
           ,x"0201" -- 235E
           ,x"c8bc" -- 2360
           ,x"0420" -- 2362
           ,x"817c" -- 2364
           ,x"0420" -- 2366
           ,x"8170" -- 2368
           ,x"c2e0" -- 236A
           ,x"ed2c" -- 236C
           ,x"045b" -- 236E
           ,x"efa8" -- 2370
           ,x"8d74" -- 2372
           ,x"c0be" -- 2374
           ,x"c802" -- 2376
           ,x"803c" -- 2378
           ,x"04e0" -- 237A
           ,x"ed3a" -- 237C
           ,x"c060" -- 237E
           ,x"8042" -- 2380
           ,x"1304" -- 2382
           ,x"04e0" -- 2384
           ,x"8042" -- 2386
           ,x"0460" -- 2388
           ,x"94f4" -- 238A
           ,x"c042" -- 238C
           ,x"c1e0" -- 238E
           ,x"ed04" -- 2390
           ,x"0202" -- 2392
           ,x"c8d4" -- 2394
           ,x"06a0" -- 2396
           ,x"8e20" -- 2398
           ,x"0281" -- 239A
           ,x"0033" -- 239C
           ,x"1203" -- 239E
           ,x"0202" -- 23A0
           ,x"cce0" -- 23A2
           ,x"1003" -- 23A4
           ,x"a041" -- 23A6
           ,x"c0a1" -- 23A8
           ,x"8e54" -- 23AA
           ,x"06a0" -- 23AC
           ,x"8e20" -- 23AE
           ,x"0202" -- 23B0
           ,x"c8bc" -- 23B2
           ,x"06a0" -- 23B4
           ,x"8e20" -- 23B6
           ,x"c020" -- 23B8
           ,x"ede4" -- 23BA
           ,x"132d" -- 23BC
           ,x"c120" -- 23BE
           ,x"ed32" -- 23C0
           ,x"1015" -- 23C2
           ,x"c0a0" -- 23C4
           ,x"ede6" -- 23C6
           ,x"0222" -- 23C8
           ,x"fffc" -- 23CA
           ,x"8802" -- 23CC
           ,x"edd2" -- 23CE
           ,x"1a06" -- 23D0
           ,x"c120" -- 23D2
           ,x"ed32" -- 23D4
           ,x"c822" -- 23D6
           ,x"fffe" -- 23D8
           ,x"ed32" -- 23DA
           ,x"1002" -- 23DC
           ,x"c120" -- 23DE
           ,x"ed32" -- 23E0
           ,x"06a0" -- 23E2
           ,x"a214" -- 23E4
           ,x"0a0d" -- 23E6
           ,x"5374" -- 23E8
           ,x"6f70" -- 23EA
           ,x"2000" -- 23EC
           ,x"0720" -- 23EE
           ,x"803c" -- 23F0
           ,x"06a0" -- 23F2
           ,x"a218" -- 23F4
           ,x"6174" -- 23F6
           ,x"2000" -- 23F8
           ,x"c820" -- 23FA
           ,x"8020" -- 23FC
           ,x"ef9e" -- 23FE
           ,x"0420" -- 2400
           ,x"b05a" -- 2402
           ,x"c060" -- 2404
           ,x"ed12" -- 2406
           ,x"1307" -- 2408
           ,x"dde0" -- 240A
           ,x"c875" -- 240C
           ,x"c820" -- 240E
           ,x"801a" -- 2410
           ,x"ef9e" -- 2412
           ,x"0420" -- 2414
           ,x"b05a" -- 2416
           ,x"0420" -- 2418
           ,x"8190" -- 241A
           ,x"0460" -- 241C
           ,x"8124" -- 241E
           ,x"ddf2" -- 2420
           ,x"15fe" -- 2422
           ,x"1102" -- 2424
           ,x"0607" -- 2426
           ,x"045b" -- 2428
           ,x"04c9" -- 242A
           ,x"d267" -- 242C
           ,x"ffff" -- 242E
           ,x"0509" -- 2430
           ,x"d9c9" -- 2432
           ,x"ffff" -- 2434
           ,x"10f8" -- 2436
           ,x"c060" -- 2438
           ,x"ede4" -- 243A
           ,x"1307" -- 243C
           ,x"c820" -- 243E
           ,x"802e" -- 2440
           ,x"ef9e" -- 2442
           ,x"0420" -- 2444
           ,x"b558" -- 2446
           ,x"0460" -- 2448
           ,x"aefc" -- 244A
           ,x"0560" -- 244C
           ,x"804a" -- 244E
           ,x"0460" -- 2450
           ,x"8124" -- 2452
           ,x"0000" -- 2454
           ,x"ccec" -- 2456
           ,x"ccf8" -- 2458
           ,x"cd0b" -- 245A
           ,x"cd1e" -- 245C
           ,x"cd33" -- 245E
           ,x"cd45" -- 2460
           ,x"cd56" -- 2462
           ,x"cd68" -- 2464
           ,x"cd7d" -- 2466
           ,x"cd96" -- 2468
           ,x"cda3" -- 246A
           ,x"cdb1" -- 246C
           ,x"cdc0" -- 246E
           ,x"cdd3" -- 2470
           ,x"cdec" -- 2472
           ,x"ce02" -- 2474
           ,x"ce20" -- 2476
           ,x"ce36" -- 2478
           ,x"ce48" -- 247A
           ,x"ce5b" -- 247C
           ,x"0000" -- 247E
           ,x"ce74" -- 2480
           ,x"ce86" -- 2482
           ,x"ce96" -- 2484
           ,x"ceae" -- 2486
           ,x"cecc" -- 2488
           ,x"cee6" -- 248A
           ,x"cefc" -- 248C
           ,x"cf0c" -- 248E
           ,x"cf23" -- 2490
           ,x"cf2e" -- 2492
           ,x"cf3a" -- 2494
           ,x"cf45" -- 2496
           ,x"cf5d" -- 2498
           ,x"cf70" -- 249A
           ,x"cf7f" -- 249C
           ,x"cf9a" -- 249E
           ,x"cfab" -- 24A0
           ,x"cfbd" -- 24A2
           ,x"cfd3" -- 24A4
           ,x"cfe5" -- 24A6
           ,x"0000" -- 24A8
           ,x"0000" -- 24AA
           ,x"0000" -- 24AC
           ,x"0000" -- 24AE
           ,x"cfff" -- 24B0
           ,x"0000" -- 24B2
           ,x"d014" -- 24B4
           ,x"c8e2" -- 24B6
           ,x"d02b" -- 24B8
           ,x"d040" -- 24BA
           ,x"020c" -- 24BC
           ,x"eea0" -- 24BE
           ,x"020b" -- 24C0
           ,x"eeb8" -- 24C2
           ,x"0420" -- 24C4
           ,x"b4e8" -- 24C6
           ,x"1001" -- 24C8
           ,x"1016" -- 24CA
           ,x"04c2" -- 24CC
           ,x"c10c" -- 24CE
           ,x"c820" -- 24D0
           ,x"8022" -- 24D2
           ,x"ef9e" -- 24D4
           ,x"0420" -- 24D6
           ,x"b558" -- 24D8
           ,x"0280" -- 24DA
           ,x"3f00" -- 24DC
           ,x"1608" -- 24DE
           ,x"0582" -- 24E0
           ,x"c80c" -- 24E2
           ,x"ef9e" -- 24E4
           ,x"05cc" -- 24E6
           ,x"0420" -- 24E8
           ,x"b558" -- 24EA
           ,x"82cc" -- 24EC
           ,x"1af5" -- 24EE
           ,x"c6c2" -- 24F0
           ,x"0404" -- 24F2
           ,x"0460" -- 24F4
           ,x"aefc" -- 24F6
           ,x"0460" -- 24F8
           ,x"97b2" -- 24FA
           ,x"05a0" -- 24FC
           ,x"ef6a" -- 24FE
           ,x"d031" -- 2500
           ,x"130a" -- 2502
           ,x"9012" -- 2504
           ,x"16fa" -- 2506
           ,x"c0c2" -- 2508
           ,x"0583" -- 250A
           ,x"c101" -- 250C
           ,x"d033" -- 250E
           ,x"1305" -- 2510
           ,x"9d00" -- 2512
           ,x"13fc" -- 2514
           ,x"10f2" -- 2516
           ,x"04e0" -- 2518
           ,x"ef6a" -- 251A
           ,x"0460" -- 251C
           ,x"b6be" -- 251E
           ,x"9c52" -- 2520
           ,x"16fc" -- 2522
           ,x"dc92" -- 2524
           ,x"13fa" -- 2526
           ,x"05a0" -- 2528
           ,x"ef6a" -- 252A
           ,x"10f9" -- 252C
           ,x"d072" -- 252E
           ,x"13f5" -- 2530
           ,x"05a0" -- 2532
           ,x"ef6a" -- 2534
           ,x"10fb" -- 2536
           ,x"c820" -- 2538
           ,x"802c" -- 253A
           ,x"ef9e" -- 253C
           ,x"0420" -- 253E
           ,x"b558" -- 2540
           ,x"101a" -- 2542
           ,x"06a0" -- 2544
           ,x"c1aa" -- 2546
           ,x"0241" -- 2548
           ,x"000f" -- 254A
           ,x"1304" -- 254C
           ,x"0281" -- 254E
           ,x"0008" -- 2550
           ,x"1501" -- 2552
           ,x"06c3" -- 2554
           ,x"0a61" -- 2556
           ,x"0221" -- 2558
           ,x"3003" -- 255A
           ,x"100a" -- 255C
           ,x"06a0" -- 255E
           ,x"c1aa" -- 2560
           ,x"0241" -- 2562
           ,x"00ff" -- 2564
           ,x"0221" -- 2566
           ,x"1d00" -- 2568
           ,x"c0c3" -- 256A
           ,x"1602" -- 256C
           ,x"0221" -- 256E
           ,x"0100" -- 2570
           ,x"c320" -- 2572
           ,x"8040" -- 2574
           ,x"0481" -- 2576
           ,x"0460" -- 2578
           ,x"aefc" -- 257A
           ,x"06a0" -- 257C
           ,x"bbd6" -- 257E
           ,x"0241" -- 2580
           ,x"000f" -- 2582
           ,x"c001" -- 2584
           ,x"0a61" -- 2586
           ,x"0221" -- 2588
           ,x"3401" -- 258A
           ,x"c320" -- 258C
           ,x"8040" -- 258E
           ,x"0481" -- 2590
           ,x"c000" -- 2592
           ,x"1304" -- 2594
           ,x"0280" -- 2596
           ,x"0008" -- 2598
           ,x"1501" -- 259A
           ,x"0981" -- 259C
           ,x"c801" -- 259E
           ,x"ef6a" -- 25A0
           ,x"0460" -- 25A2
           ,x"b6be" -- 25A4
           ,x"06a0" -- 25A6
           ,x"bbd6" -- 25A8
           ,x"0241" -- 25AA
           ,x"00ff" -- 25AC
           ,x"0221" -- 25AE
           ,x"1f00" -- 25B0
           ,x"c320" -- 25B2
           ,x"8040" -- 25B4
           ,x"0481" -- 25B6
           ,x"16f4" -- 25B8
           ,x"05a0" -- 25BA
           ,x"ef6a" -- 25BC
           ,x"10f1" -- 25BE
           ,x"c020" -- 25C0
           ,x"ede4" -- 25C2
           ,x"130d" -- 25C4
           ,x"04c0" -- 25C6
           ,x"d038" -- 25C8
           ,x"0701" -- 25CA
           ,x"0581" -- 25CC
           ,x"9838" -- 25CE
           ,x"ab26" -- 25D0
           ,x"16fc" -- 25D2
           ,x"c0e0" -- 25D4
           ,x"ed0c" -- 25D6
           ,x"0960" -- 25D8
           ,x"a0c0" -- 25DA
           ,x"ccc8" -- 25DC
           ,x"c4c1" -- 25DE
           ,x"0460" -- 25E0
           ,x"af02" -- 25E2
           ,x"04c0" -- 25E4
           ,x"d038" -- 25E6
           ,x"0280" -- 25E8
           ,x"4300" -- 25EA
           ,x"1601" -- 25EC
           ,x"d038" -- 25EE
           ,x"0280" -- 25F0
           ,x"7400" -- 25F2
           ,x"1a59" -- 25F4
           ,x"c3a0" -- 25F6
           ,x"edd6" -- 25F8
           ,x"0970" -- 25FA
           ,x"a380" -- 25FC
           ,x"022e" -- 25FE
           ,x"ff20" -- 2600
           ,x"c05e" -- 2602
           ,x"161e" -- 2604
           ,x"0705" -- 2606
           ,x"06a0" -- 2608
           ,x"b6d4" -- 260A
           ,x"04f6" -- 260C
           ,x"1002" -- 260E
           ,x"06a0" -- 2610
           ,x"b6dc" -- 2612
           ,x"06a0" -- 2614
           ,x"bbd6" -- 2616
           ,x"0646" -- 2618
           ,x"c0d6" -- 261A
           ,x"0583" -- 261C
           ,x"cd81" -- 261E
           ,x"0736" -- 2620
           ,x"cd83" -- 2622
           ,x"0280" -- 2624
           ,x"3f00" -- 2626
           ,x"13f3" -- 2628
           ,x"0280" -- 262A
           ,x"4b00" -- 262C
           ,x"1607" -- 262E
           ,x"0646" -- 2630
           ,x"c016" -- 2632
           ,x"c280" -- 2634
           ,x"0a2a" -- 2636
           ,x"0201" -- 2638
           ,x"0001" -- 263A
           ,x"1011" -- 263C
           ,x"0460" -- 263E
           ,x"aef2" -- 2640
           ,x"0608" -- 2642
           ,x"0420" -- 2644
           ,x"b526" -- 2646
           ,x"1026" -- 2648
           ,x"0226" -- 264A
           ,x"fffc" -- 264C
           ,x"c096" -- 264E
           ,x"0582" -- 2650
           ,x"3881" -- 2652
           ,x"c082" -- 2654
           ,x"1626" -- 2656
           ,x"c043" -- 2658
           ,x"1124" -- 265A
           ,x"c981" -- 265C
           ,x"fffe" -- 265E
           ,x"0600" -- 2660
           ,x"16f3" -- 2662
           ,x"0226" -- 2664
           ,x"fffc" -- 2666
           ,x"c016" -- 2668
           ,x"0580" -- 266A
           ,x"3840" -- 266C
           ,x"38a0" -- 266E
           ,x"b92a" -- 2670
           ,x"c082" -- 2672
           ,x"1617" -- 2674
           ,x"a0ca" -- 2676
           ,x"c0a0" -- 2678
           ,x"edda" -- 267A
           ,x"6083" -- 267C
           ,x"8802" -- 267E
           ,x"edd8" -- 2680
           ,x"1a10" -- 2682
           ,x"c782" -- 2684
           ,x"c802" -- 2686
           ,x"edda" -- 2688
           ,x"ccb6" -- 268A
           ,x"05a6" -- 268C
           ,x"fffe" -- 268E
           ,x"16fc" -- 2690
           ,x"04c0" -- 2692
           ,x"d038" -- 2694
           ,x"0280" -- 2696
           ,x"3f00" -- 2698
           ,x"13a4" -- 269A
           ,x"c800" -- 269C
           ,x"ede8" -- 269E
           ,x"0460" -- 26A0
           ,x"aefc" -- 26A2
           ,x"0460" -- 26A4
           ,x"a5a6" -- 26A6
           ,x"0420" -- 26A8
           ,x"8d70" -- 26AA
           ,x"0010" -- 26AC
           ,x"0420" -- 26AE
           ,x"b4e8" -- 26B0
           ,x"1003" -- 26B2
           ,x"1002" -- 26B4
           ,x"0460" -- 26B6
           ,x"9844" -- 26B8
           ,x"c1e0" -- 26BA
           ,x"ed04" -- 26BC
           ,x"0205" -- 26BE
           ,x"0084" -- 26C0
           ,x"ddf2" -- 26C2
           ,x"1304" -- 26C4
           ,x"0605" -- 26C6
           ,x"16fc" -- 26C8
           ,x"0460" -- 26CA
           ,x"93fc" -- 26CC
           ,x"c160" -- 26CE
           ,x"ede6" -- 26D0
           ,x"c825" -- 26D2
           ,x"fffe" -- 26D4
           ,x"ed32" -- 26D6
           ,x"06a0" -- 26D8
           ,x"a374" -- 26DA
           ,x"4820" -- 26DC
           ,x"b920" -- 26DE
           ,x"8046" -- 26E0
           ,x"c060" -- 26E2
           ,x"ed32" -- 26E4
           ,x"06a0" -- 26E6
           ,x"a2a6" -- 26E8
           ,x"c808" -- 26EA
           ,x"ede6" -- 26EC
           ,x"0460" -- 26EE
           ,x"af02" -- 26F0
           ,x"04e0" -- 26F2
           ,x"8046" -- 26F4
           ,x"1002" -- 26F6
           ,x"0720" -- 26F8
           ,x"8046" -- 26FA
           ,x"0460" -- 26FC
           ,x"aef8" -- 26FE
           ,x"06a0" -- 2700
           ,x"9284" -- 2702
           ,x"c0d4" -- 2704
           ,x"160a" -- 2706
           ,x"c0e0" -- 2708
           ,x"edda" -- 270A
           ,x"0223" -- 270C
           ,x"fffa" -- 270E
           ,x"8803" -- 2710
           ,x"edd8" -- 2712
           ,x"1a70" -- 2714
           ,x"c503" -- 2716
           ,x"c803" -- 2718
           ,x"edda" -- 271A
           ,x"c120" -- 271C
           ,x"ed08" -- 271E
           ,x"9838" -- 2720
           ,x"ab26" -- 2722
           ,x"1664" -- 2724
           ,x"c014" -- 2726
           ,x"1315" -- 2728
           ,x"8001" -- 272A
           ,x"1307" -- 272C
           ,x"0224" -- 272E
           ,x"0012" -- 2730
           ,x"8804" -- 2732
           ,x"ed06" -- 2734
           ,x"1af7" -- 2736
           ,x"0460" -- 2738
           ,x"9576" -- 273A
           ,x"06a0" -- 273C
           ,x"9142" -- 273E
           ,x"10f2" -- 2740
           ,x"c144" -- 2742
           ,x"c004" -- 2744
           ,x"0220" -- 2746
           ,x"0012" -- 2748
           ,x"cd70" -- 274A
           ,x"8800" -- 274C
           ,x"ed06" -- 274E
           ,x"12fc" -- 2750
           ,x"045b" -- 2752
           ,x"cd01" -- 2754
           ,x"0420" -- 2756
           ,x"b540" -- 2758
           ,x"0280" -- 275A
           ,x"3800" -- 275C
           ,x"1649" -- 275E
           ,x"c183" -- 2760
           ,x"ccf2" -- 2762
           ,x"ccf2" -- 2764
           ,x"c4d2" -- 2766
           ,x"04f4" -- 2768
           ,x"04d4" -- 276A
           ,x"05b4" -- 276C
           ,x"04f4" -- 276E
           ,x"0420" -- 2770
           ,x"b540" -- 2772
           ,x"c1c4" -- 2774
           ,x"cd32" -- 2776
           ,x"cd32" -- 2778
           ,x"cd12" -- 277A
           ,x"04c5" -- 277C
           ,x"0280" -- 277E
           ,x"3a00" -- 2780
           ,x"160c" -- 2782
           ,x"0420" -- 2784
           ,x"b540" -- 2786
           ,x"c044" -- 2788
           ,x"0221" -- 278A
           ,x"fff4" -- 278C
           ,x"c152" -- 278E
           ,x"1602" -- 2790
           ,x"c162" -- 2792
           ,x"0002" -- 2794
           ,x"cc72" -- 2796
           ,x"cc72" -- 2798
           ,x"c452" -- 279A
           ,x"c508" -- 279C
           ,x"0634" -- 279E
           ,x"c520" -- 27A0
           ,x"ede6" -- 27A2
           ,x"c086" -- 27A4
           ,x"c047" -- 27A6
           ,x"06a0" -- 27A8
           ,x"b9be" -- 27AA
           ,x"c072" -- 27AC
           ,x"1602" -- 27AE
           ,x"c052" -- 27B0
           ,x"131b" -- 27B2
           ,x"2845" -- 27B4
           ,x"1119" -- 27B6
           ,x"c164" -- 27B8
           ,x"fff0" -- 27BA
           ,x"04e4" -- 27BC
           ,x"fff0" -- 27BE
           ,x"c1a0" -- 27C0
           ,x"ede6" -- 27C2
           ,x"0226" -- 27C4
           ,x"fffc" -- 27C6
           ,x"8806" -- 27C8
           ,x"edd2" -- 27CA
           ,x"1a16" -- 27CC
           ,x"c216" -- 27CE
           ,x"a220" -- 27D0
           ,x"ed0e" -- 27D2
           ,x"9838" -- 27D4
           ,x"ab81" -- 27D6
           ,x"16f5" -- 27D8
           ,x"06a0" -- 27DA
           ,x"9284" -- 27DC
           ,x"8141" -- 27DE
           ,x"16f1" -- 27E0
           ,x"c806" -- 27E2
           ,x"ede6" -- 27E4
           ,x"0460" -- 27E6
           ,x"aef8" -- 27E8
           ,x"0460" -- 27EA
           ,x"aefc" -- 27EC
           ,x"0460" -- 27EE
           ,x"9802" -- 27F0
           ,x"0460" -- 27F2
           ,x"aef2" -- 27F4
           ,x"0460" -- 27F6
           ,x"a5a6" -- 27F8
           ,x"0420" -- 27FA
           ,x"8d70" -- 27FC
           ,x"001f" -- 27FE
           ,x"0420" -- 2800
           ,x"8d70" -- 2802
           ,x"0014" -- 2804
           ,x"06a0" -- 2806
           ,x"9284" -- 2808
           ,x"c194" -- 280A
           ,x"1309" -- 280C
           ,x"c120" -- 280E
           ,x"ed08" -- 2810
           ,x"8d01" -- 2812
           ,x"1308" -- 2814
           ,x"0224" -- 2816
           ,x"0010" -- 2818
           ,x"8804" -- 281A
           ,x"ed06" -- 281C
           ,x"1af9" -- 281E
           ,x"0420" -- 2820
           ,x"8d70" -- 2822
           ,x"0020" -- 2824
           ,x"c084" -- 2826
           ,x"c172" -- 2828
           ,x"160f" -- 282A
           ,x"c152" -- 282C
           ,x"c2c6" -- 282E
           ,x"c07b" -- 2830
           ,x"160b" -- 2832
           ,x"c064" -- 2834
           ,x"0006" -- 2836
           ,x"1608" -- 2838
           ,x"c05b" -- 283A
           ,x"a052" -- 283C
           ,x"1901" -- 283E
           ,x"1004" -- 2840
           ,x"c6c1" -- 2842
           ,x"6064" -- 2844
           ,x"0008" -- 2846
           ,x"1010" -- 2848
           ,x"c046" -- 284A
           ,x"c084" -- 284C
           ,x"06a0" -- 284E
           ,x"b98e" -- 2850
           ,x"c042" -- 2852
           ,x"cdb1" -- 2854
           ,x"cdb1" -- 2856
           ,x"c591" -- 2858
           ,x"c044" -- 285A
           ,x"0221" -- 285C
           ,x"0006" -- 285E
           ,x"06a0" -- 2860
           ,x"b9be" -- 2862
           ,x"c072" -- 2864
           ,x"1602" -- 2866
           ,x"c052" -- 2868
           ,x"1305" -- 286A
           ,x"2845" -- 286C
           ,x"1103" -- 286E
           ,x"04e4" -- 2870
           ,x"fffe" -- 2872
           ,x"1005" -- 2874
           ,x"c224" -- 2876
           ,x"000c" -- 2878
           ,x"c824" -- 287A
           ,x"000e" -- 287C
           ,x"ede6" -- 287E
           ,x"0460" -- 2880
           ,x"aef8" -- 2882
           ,x"04c0" -- 2884
           ,x"d038" -- 2886
           ,x"0280" -- 2888
           ,x"7400" -- 288A
           ,x"1ab9" -- 288C
           ,x"c120" -- 288E
           ,x"edd4" -- 2890
           ,x"0970" -- 2892
           ,x"a100" -- 2894
           ,x"c064" -- 2896
           ,x"ff20" -- 2898
           ,x"11b2" -- 289A
           ,x"c120" -- 289C
           ,x"edd6" -- 289E
           ,x"a100" -- 28A0
           ,x"0224" -- 28A2
           ,x"ff20" -- 28A4
           ,x"045b" -- 28A6
           ,x"c209" -- 28A8
           ,x"c187" -- 28AA
           ,x"04c3" -- 28AC
           ,x"04c4" -- 28AE
           ,x"04c5" -- 28B0
           ,x"06a0" -- 28B2
           ,x"9396" -- 28B4
           ,x"100a" -- 28B6
           ,x"1002" -- 28B8
           ,x"0703" -- 28BA
           ,x"1004" -- 28BC
           ,x"c0c3" -- 28BE
           ,x"1601" -- 28C0
           ,x"0584" -- 28C2
           ,x"0585" -- 28C4
           ,x"dda0" -- 28C6
           ,x"c8d6" -- 28C8
           ,x"10f3" -- 28CA
           ,x"022a" -- 28CC
           ,x"fff3" -- 28CE
           ,x"050a" -- 28D0
           ,x"810a" -- 28D2
           ,x"151a" -- 28D4
           ,x"6144" -- 28D6
           ,x"a14a" -- 28D8
           ,x"0285" -- 28DA
           ,x"000c" -- 28DC
           ,x"1102" -- 28DE
           ,x"0205" -- 28E0
           ,x"000c" -- 28E2
           ,x"c005" -- 28E4
           ,x"0600" -- 28E6
           ,x"06a0" -- 28E8
           ,x"b1e8" -- 28EA
           ,x"058a" -- 28EC
           ,x"c209" -- 28EE
           ,x"04c5" -- 28F0
           ,x"06a0" -- 28F2
           ,x"9396" -- 28F4
           ,x"100a" -- 28F6
           ,x"100c" -- 28F8
           ,x"102c" -- 28FA
           ,x"0280" -- 28FC
           ,x"2c00" -- 28FE
           ,x"1602" -- 2900
           ,x"c145" -- 2902
           ,x"1320" -- 2904
           ,x"ddc0" -- 2906
           ,x"10f4" -- 2908
           ,x"c1c6" -- 290A
           ,x"cb47" -- 290C
           ,x"000e" -- 290E
           ,x"0380" -- 2910
           ,x"0604" -- 2912
           ,x"8284" -- 2914
           ,x"111b" -- 2916
           ,x"1302" -- 2918
           ,x"c104" -- 291A
           ,x"1611" -- 291C
           ,x"0280" -- 291E
           ,x"2400" -- 2920
           ,x"13f1" -- 2922
           ,x"0280" -- 2924
           ,x"5300" -- 2926
           ,x"1605" -- 2928
           ,x"c30c" -- 292A
           ,x"130c" -- 292C
           ,x"0200" -- 292E
           ,x"2d00" -- 2930
           ,x"10e9" -- 2932
           ,x"0280" -- 2934
           ,x"3c00" -- 2936
           ,x"1603" -- 2938
           ,x"c30c" -- 293A
           ,x"16e4" -- 293C
           ,x"1003" -- 293E
           ,x"0280" -- 2940
           ,x"3000" -- 2942
           ,x"1302" -- 2944
           ,x"0200" -- 2946
           ,x"2000" -- 2948
           ,x"ddc0" -- 294A
           ,x"10d2" -- 294C
           ,x"06a0" -- 294E
           ,x"9384" -- 2950
           ,x"10cf" -- 2952
           ,x"ddc0" -- 2954
           ,x"06a0" -- 2956
           ,x"9396" -- 2958
           ,x"10cd" -- 295A
           ,x"100a" -- 295C
           ,x"1000" -- 295E
           ,x"0280" -- 2960
           ,x"3e00" -- 2962
           ,x"1604" -- 2964
           ,x"c30c" -- 2966
           ,x"1602" -- 2968
           ,x"0200" -- 296A
           ,x"2000" -- 296C
           ,x"ddc0" -- 296E
           ,x"10f2" -- 2970
           ,x"0604" -- 2972
           ,x"8284" -- 2974
           ,x"1103" -- 2976
           ,x"0200" -- 2978
           ,x"3000" -- 297A
           ,x"10f8" -- 297C
           ,x"06a0" -- 297E
           ,x"9384" -- 2980
           ,x"10e9" -- 2982
           ,x"060a" -- 2984
           ,x"0705" -- 2986
           ,x"ddf3" -- 2988
           ,x"1604" -- 298A
           ,x"0607" -- 298C
           ,x"0603" -- 298E
           ,x"dde0" -- 2990
           ,x"b0f7" -- 2992
           ,x"045b" -- 2994
           ,x"04c0" -- 2996
           ,x"d038" -- 2998
           ,x"1323" -- 299A
           ,x"0280" -- 299C
           ,x"3c00" -- 299E
           ,x"131f" -- 29A0
           ,x"0280" -- 29A2
           ,x"2400" -- 29A4
           ,x"131c" -- 29A6
           ,x"0280" -- 29A8
           ,x"5300" -- 29AA
           ,x"1319" -- 29AC
           ,x"0280" -- 29AE
           ,x"3000" -- 29B0
           ,x"1316" -- 29B2
           ,x"0280" -- 29B4
           ,x"3900" -- 29B6
           ,x"1313" -- 29B8
           ,x"0280" -- 29BA
           ,x"2e00" -- 29BC
           ,x"130f" -- 29BE
           ,x"0280" -- 29C0
           ,x"4500" -- 29C2
           ,x"1606" -- 29C4
           ,x"0200" -- 29C6
           ,x"2000" -- 29C8
           ,x"c30c" -- 29CA
           ,x"1302" -- 29CC
           ,x"0200" -- 29CE
           ,x"2d00" -- 29D0
           ,x"0280" -- 29D2
           ,x"5e00" -- 29D4
           ,x"1602" -- 29D6
           ,x"0200" -- 29D8
           ,x"2e00" -- 29DA
           ,x"05cb" -- 29DC
           ,x"05cb" -- 29DE
           ,x"05cb" -- 29E0
           ,x"045b" -- 29E2
           ,x"06a0" -- 29E4
           ,x"bbd6" -- 29E6
           ,x"0281" -- 29E8
           ,x"000b" -- 29EA
           ,x"1604" -- 29EC
           ,x"d060" -- 29EE
           ,x"0000" -- 29F0
           ,x"0981" -- 29F2
           ,x"101d" -- 29F4
           ,x"0281" -- 29F6
           ,x"0014" -- 29F8
           ,x"1203" -- 29FA
           ,x"0420" -- 29FC
           ,x"8d70" -- 29FE
           ,x"0023" -- 2A00
           ,x"a041" -- 2A02
           ,x"c061" -- 2A04
           ,x"803a" -- 2A06
           ,x"1013" -- 2A08
           ,x"c052" -- 2A0A
           ,x"1317" -- 2A0C
           ,x"c802" -- 2A0E
           ,x"ef7e" -- 2A10
           ,x"0420" -- 2A12
           ,x"bc3e" -- 2A14
           ,x"0241" -- 2A16
           ,x"7f00" -- 2A18
           ,x"8801" -- 2A1A
           ,x"c838" -- 2A1C
           ,x"140c" -- 2A1E
           ,x"c820" -- 2A20
           ,x"c83a" -- 2A22
           ,x"ef7e" -- 2A24
           ,x"0420" -- 2A26
           ,x"bf7c" -- 2A28
           ,x"0420" -- 2A2A
           ,x"bd46" -- 2A2C
           ,x"1004" -- 2A2E
           ,x"0420" -- 2A30
           ,x"be74" -- 2A32
           ,x"c801" -- 2A34
           ,x"ef6a" -- 2A36
           ,x"0202" -- 2A38
           ,x"ef68" -- 2A3A
           ,x"0460" -- 2A3C
           ,x"b6ac" -- 2A3E
           ,x"c802" -- 2A40
           ,x"ef7e" -- 2A42
           ,x"0420" -- 2A44
           ,x"bc3e" -- 2A46
           ,x"c052" -- 2A48
           ,x"1304" -- 2A4A
           ,x"15f7" -- 2A4C
           ,x"0420" -- 2A4E
           ,x"bd0c" -- 2A50
           ,x"10f2" -- 2A52
           ,x"0760" -- 2A54
           ,x"ef6a" -- 2A56
           ,x"19ef" -- 2A58
           ,x"0200" -- 2A5A
           ,x"4480" -- 2A5C
           ,x"04c2" -- 2A5E
           ,x"c820" -- 2A60
           ,x"8016" -- 2A62
           ,x"ef7e" -- 2A64
           ,x"0420" -- 2A66
           ,x"bc3e" -- 2A68
           ,x"10e6" -- 2A6A
           ,x"0420" -- 2A6C
           ,x"8194" -- 2A6E
           ,x"10e3" -- 2A70
           ,x"1000" -- 2A72
           ,x"06c0" -- 2A74
           ,x"06a0" -- 2A76
           ,x"bbd6" -- 2A78
           ,x"c041" -- 2A7A
           ,x"1302" -- 2A7C
           ,x"8040" -- 2A7E
           ,x"16db" -- 2A80
           ,x"c040" -- 2A82
           ,x"10d5" -- 2A84
           ,x"c012" -- 2A86
           ,x"1603" -- 2A88
           ,x"0202" -- 2A8A
           ,x"ef68" -- 2A8C
           ,x"045b" -- 2A8E
           ,x"0240" -- 2A90
           ,x"7f00" -- 2A92
           ,x"0280" -- 2A94
           ,x"4900" -- 2A96
           ,x"15f8" -- 2A98
           ,x"c802" -- 2A9A
           ,x"ef7e" -- 2A9C
           ,x"0420" -- 2A9E
           ,x"bc3e" -- 2AA0
           ,x"0280" -- 2AA2
           ,x"4100" -- 2AA4
           ,x"11f1" -- 2AA6
           ,x"c820" -- 2AA8
           ,x"8012" -- 2AAA
           ,x"ef7e" -- 2AAC
           ,x"0420" -- 2AAE
           ,x"bc32" -- 2AB0
           ,x"c820" -- 2AB2
           ,x"c83a" -- 2AB4
           ,x"ef7e" -- 2AB6
           ,x"0420" -- 2AB8
           ,x"bf7c" -- 2ABA
           ,x"0420" -- 2ABC
           ,x"bd46" -- 2ABE
           ,x"0420" -- 2AC0
           ,x"bd0c" -- 2AC2
           ,x"c820" -- 2AC4
           ,x"8012" -- 2AC6
           ,x"ef7e" -- 2AC8
           ,x"0420" -- 2ACA
           ,x"bc4a" -- 2ACC
           ,x"10dd" -- 2ACE
           ,x"c0c1" -- 2AD0
           ,x"1502" -- 2AD2
           ,x"0460" -- 2AD4
           ,x"bc10" -- 2AD6
           ,x"06a0" -- 2AD8
           ,x"bbd6" -- 2ADA
           ,x"c281" -- 2ADC
           ,x"0741" -- 2ADE
           ,x"04c0" -- 2AE0
           ,x"3c03" -- 2AE2
           ,x"c28a" -- 2AE4
           ,x"15a4" -- 2AE6
           ,x"13a3" -- 2AE8
           ,x"c041" -- 2AEA
           ,x"13a1" -- 2AEC
           ,x"0501" -- 2AEE
           ,x"a043" -- 2AF0
           ,x"109e" -- 2AF2
           ,x"c160" -- 2AF4
           ,x"ede6" -- 2AF6
           ,x"c825" -- 2AF8
           ,x"fffe" -- 2AFA
           ,x"803e" -- 2AFC
           ,x"04c6" -- 2AFE
           ,x"102a" -- 2B00
           ,x"c160" -- 2B02
           ,x"ede6" -- 2B04
           ,x"1031" -- 2B06
           ,x"c160" -- 2B08
           ,x"ede6" -- 2B0A
           ,x"1024" -- 2B0C
           ,x"04c3" -- 2B0E
           ,x"1001" -- 2B10
           ,x"0703" -- 2B12
           ,x"c188" -- 2B14
           ,x"05c6" -- 2B16
           ,x"04c0" -- 2B18
           ,x"d036" -- 2B1A
           ,x"1306" -- 2B1C
           ,x"0280" -- 2B1E
           ,x"3c00" -- 2B20
           ,x"1313" -- 2B22
           ,x"0280" -- 2B24
           ,x"4700" -- 2B26
           ,x"162c" -- 2B28
           ,x"c160" -- 2B2A
           ,x"ede6" -- 2B2C
           ,x"130d" -- 2B2E
           ,x"c0c3" -- 2B30
           ,x"130b" -- 2B32
           ,x"c185" -- 2B34
           ,x"0226" -- 2B36
           ,x"fffc" -- 2B38
           ,x"8806" -- 2B3A
           ,x"edd2" -- 2B3C
           ,x"1a19" -- 2B3E
           ,x"c806" -- 2B40
           ,x"ede6" -- 2B42
           ,x"c196" -- 2B44
           ,x"a1a0" -- 2B46
           ,x"ed0e" -- 2B48
           ,x"d078" -- 2B4A
           ,x"06c1" -- 2B4C
           ,x"d078" -- 2B4E
           ,x"06c1" -- 2B50
           ,x"0922" -- 2B52
           ,x"130a" -- 2B54
           ,x"c0e0" -- 2B56
           ,x"eddc" -- 2B58
           ,x"8803" -- 2B5A
           ,x"ed08" -- 2B5C
           ,x"140b" -- 2B5E
           ,x"ccc6" -- 2B60
           ,x"cce0" -- 2B62
           ,x"ede6" -- 2B64
           ,x"c803" -- 2B66
           ,x"eddc" -- 2B68
           ,x"06a0" -- 2B6A
           ,x"a2a6" -- 2B6C
           ,x"0460" -- 2B6E
           ,x"af24" -- 2B70
           ,x"04c6" -- 2B72
           ,x"10ea" -- 2B74
           ,x"0420" -- 2B76
           ,x"8d70" -- 2B78
           ,x"000b" -- 2B7A
           ,x"0420" -- 2B7C
           ,x"8d70" -- 2B7E
           ,x"000c" -- 2B80
           ,x"0420" -- 2B82
           ,x"8d70" -- 2B84
           ,x"0025" -- 2B86
           ,x"c0e0" -- 2B88
           ,x"eddc" -- 2B8A
           ,x"8803" -- 2B8C
           ,x"ed0a" -- 2B8E
           ,x"12f5" -- 2B90
           ,x"0643" -- 2B92
           ,x"c153" -- 2B94
           ,x"0643" -- 2B96
           ,x"c803" -- 2B98
           ,x"eddc" -- 2B9A
           ,x"c805" -- 2B9C
           ,x"ede6" -- 2B9E
           ,x"1309" -- 2BA0
           ,x"c825" -- 2BA2
           ,x"fffe" -- 2BA4
           ,x"ed32" -- 2BA6
           ,x"c213" -- 2BA8
           ,x"1302" -- 2BAA
           ,x"0460" -- 2BAC
           ,x"af38" -- 2BAE
           ,x"0460" -- 2BB0
           ,x"af16" -- 2BB2
           ,x"0460" -- 2BB4
           ,x"8124" -- 2BB6
           ,x"8820" -- 2BB8
           ,x"eddc" -- 2BBA
           ,x"ed0a" -- 2BBC
           ,x"12de" -- 2BBE
           ,x"6820" -- 2BC0
           ,x"b922" -- 2BC2
           ,x"eddc" -- 2BC4
           ,x"0460" -- 2BC6
           ,x"aef8" -- 2BC8
           ,x"04e0" -- 2BCA
           ,x"ed38" -- 2BCC
           ,x"0420" -- 2BCE
           ,x"b4e8" -- 2BD0
           ,x"1008" -- 2BD2
           ,x"1007" -- 2BD4
           ,x"0420" -- 2BD6
           ,x"b540" -- 2BD8
           ,x"c072" -- 2BDA
           ,x"161b" -- 2BDC
           ,x"c052" -- 2BDE
           ,x"1619" -- 2BE0
           ,x"1034" -- 2BE2
           ,x"0280" -- 2BE4
           ,x"3b00" -- 2BE6
           ,x"1603" -- 2BE8
           ,x"d052" -- 2BEA
           ,x"1613" -- 2BEC
           ,x"102e" -- 2BEE
           ,x"06c0" -- 2BF0
           ,x"0220" -- 2BF2
           ,x"ffab" -- 2BF4
           ,x"1502" -- 2BF6
           ,x"0460" -- 2BF8
           ,x"aef2" -- 2BFA
           ,x"0280" -- 2BFC
           ,x"0006" -- 2BFE
           ,x"15fb" -- 2C00
           ,x"c180" -- 2C02
           ,x"c0c2" -- 2C04
           ,x"0705" -- 2C06
           ,x"0420" -- 2C08
           ,x"b4e8" -- 2C0A
           ,x"100c" -- 2C0C
           ,x"100b" -- 2C0E
           ,x"0460" -- 2C10
           ,x"9844" -- 2C12
           ,x"0460" -- 2C14
           ,x"aefc" -- 2C16
           ,x"d072" -- 2C18
           ,x"1601" -- 2C1A
           ,x"0701" -- 2C1C
           ,x"7044" -- 2C1E
           ,x"160f" -- 2C20
           ,x"0605" -- 2C22
           ,x"130f" -- 2C24
           ,x"0280" -- 2C26
           ,x"3f00" -- 2C28
           ,x"1605" -- 2C2A
           ,x"c820" -- 2C2C
           ,x"8022" -- 2C2E
           ,x"ef9e" -- 2C30
           ,x"0420" -- 2C32
           ,x"b558" -- 2C34
           ,x"0200" -- 2C36
           ,x"0004" -- 2C38
           ,x"d133" -- 2C3A
           ,x"16ed" -- 2C3C
           ,x"d072" -- 2C3E
           ,x"1503" -- 2C40
           ,x"1601" -- 2C42
           ,x"0600" -- 2C44
           ,x"0640" -- 2C46
           ,x"2180" -- 2C48
           ,x"13e4" -- 2C4A
           ,x"0720" -- 2C4C
           ,x"ed38" -- 2C4E
           ,x"0460" -- 2C50
           ,x"af02" -- 2C52
           ,x"04e0" -- 2C54
           ,x"803a" -- 2C56
           ,x"04e0" -- 2C58
           ,x"ed3c" -- 2C5A
           ,x"1006" -- 2C5C
           ,x"c820" -- 2C5E
           ,x"8010" -- 2C60
           ,x"ef9e" -- 2C62
           ,x"0420" -- 2C64
           ,x"b558" -- 2C66
           ,x"0608" -- 2C68
           ,x"070f" -- 2C6A
           ,x"058f" -- 2C6C
           ,x"06a0" -- 2C6E
           ,x"8724" -- 2C70
           ,x"5400" -- 2C72
           ,x"543c" -- 2C74
           ,x"5447" -- 2C76
           ,x"fc3f" -- 2C78
           ,x"fd40" -- 2C7A
           ,x"343e" -- 2C7C
           ,x"f641" -- 2C7E
           ,x"3242" -- 2C80
           ,x"0000" -- 2C82
           ,x"0608" -- 2C84
           ,x"0420" -- 2C86
           ,x"b4e8" -- 2C88
           ,x"102d" -- 2C8A
           ,x"1039" -- 2C8C
           ,x"0420" -- 2C8E
           ,x"b526" -- 2C90
           ,x"c182" -- 2C92
           ,x"0202" -- 2C94
           ,x"c8da" -- 2C96
           ,x"06a0" -- 2C98
           ,x"971e" -- 2C9A
           ,x"0420" -- 2C9C
           ,x"b288" -- 2C9E
           ,x"100c" -- 2CA0
           ,x"04c1" -- 2CA2
           ,x"1000" -- 2CA4
           ,x"c000" -- 2CA6
           ,x"160f" -- 2CA8
           ,x"04f6" -- 2CAA
           ,x"cd81" -- 2CAC
           ,x"04f6" -- 2CAE
           ,x"04e0" -- 2CB0
           ,x"ed3c" -- 2CB2
           ,x"04e0" -- 2CB4
           ,x"ed3a" -- 2CB6
           ,x"10d7" -- 2CB8
           ,x"c000" -- 2CBA
           ,x"1605" -- 2CBC
           ,x"c806" -- 2CBE
           ,x"ef7e" -- 2CC0
           ,x"0420" -- 2CC2
           ,x"bc32" -- 2CC4
           ,x"10f4" -- 2CC6
           ,x"0202" -- 2CC8
           ,x"c8d9" -- 2CCA
           ,x"c060" -- 2CCC
           ,x"803a" -- 2CCE
           ,x"13e3" -- 2CD0
           ,x"0700" -- 2CD2
           ,x"1046" -- 2CD4
           ,x"0720" -- 2CD6
           ,x"ed3c" -- 2CD8
           ,x"c820" -- 2CDA
           ,x"800e" -- 2CDC
           ,x"ef9e" -- 2CDE
           ,x"0420" -- 2CE0
           ,x"b558" -- 2CE2
           ,x"10c1" -- 2CE4
           ,x"020b" -- 2CE6
           ,x"9668" -- 2CE8
           ,x"c34b" -- 2CEA
           ,x"c1e0" -- 2CEC
           ,x"ed04" -- 2CEE
           ,x"0205" -- 2CF0
           ,x"0084" -- 2CF2
           ,x"06a0" -- 2CF4
           ,x"99ba" -- 2CF6
           ,x"1000" -- 2CF8
           ,x"c2cd" -- 2CFA
           ,x"0460" -- 2CFC
           ,x"9772" -- 2CFE
           ,x"c182" -- 2D00
           ,x"0202" -- 2D02
           ,x"c8dd" -- 2D04
           ,x"06a0" -- 2D06
           ,x"971e" -- 2D08
           ,x"c087" -- 2D0A
           ,x"c1c6" -- 2D0C
           ,x"0205" -- 2D0E
           ,x"0064" -- 2D10
           ,x"06a0" -- 2D12
           ,x"99ba" -- 2D14
           ,x"10cc" -- 2D16
           ,x"10cb" -- 2D18
           ,x"0460" -- 2D1A
           ,x"9782" -- 2D1C
           ,x"c38b" -- 2D1E
           ,x"c3cf" -- 2D20
           ,x"1602" -- 2D22
           ,x"06a0" -- 2D24
           ,x"96ea" -- 2D26
           ,x"c1e0" -- 2D28
           ,x"ed04" -- 2D2A
           ,x"c120" -- 2D2C
           ,x"ed3a" -- 2D2E
           ,x"1602" -- 2D30
           ,x"0204" -- 2D32
           ,x"0080" -- 2D34
           ,x"0420" -- 2D36
           ,x"8198" -- 2D38
           ,x"06a0" -- 2D3A
           ,x"9d3a" -- 2D3C
           ,x"1006" -- 2D3E
           ,x"100c" -- 2D40
           ,x"0420" -- 2D42
           ,x"816c" -- 2D44
           ,x"0604" -- 2D46
           ,x"16f6" -- 2D48
           ,x"1003" -- 2D4A
           ,x"c020" -- 2D4C
           ,x"ed3c" -- 2D4E
           ,x"16f2" -- 2D50
           ,x"75d7" -- 2D52
           ,x"c1e0" -- 2D54
           ,x"ed04" -- 2D56
           ,x"045e" -- 2D58
           ,x"c060" -- 2D5A
           ,x"803a" -- 2D5C
           ,x"13eb" -- 2D5E
           ,x"06c0" -- 2D60
           ,x"c800" -- 2D62
           ,x"803a" -- 2D64
           ,x"04e0" -- 2D66
           ,x"ed3a" -- 2D68
           ,x"04e0" -- 2D6A
           ,x"ed3c" -- 2D6C
           ,x"0460" -- 2D6E
           ,x"94f4" -- 2D70
           ,x"c34b" -- 2D72
           ,x"06a0" -- 2D74
           ,x"9792" -- 2D76
           ,x"c1e0" -- 2D78
           ,x"ed04" -- 2D7A
           ,x"045d" -- 2D7C
           ,x"06a0" -- 2D7E
           ,x"9792" -- 2D80
           ,x"04e0" -- 2D82
           ,x"ed3a" -- 2D84
           ,x"c3cf" -- 2D86
           ,x"1602" -- 2D88
           ,x"0420" -- 2D8A
           ,x"8170" -- 2D8C
           ,x"0460" -- 2D8E
           ,x"aefc" -- 2D90
           ,x"8807" -- 2D92
           ,x"ed04" -- 2D94
           ,x"1302" -- 2D96
           ,x"0420" -- 2D98
           ,x"8190" -- 2D9A
           ,x"c020" -- 2D9C
           ,x"ed34" -- 2D9E
           ,x"a007" -- 2DA0
           ,x"6020" -- 2DA2
           ,x"ed04" -- 2DA4
           ,x"0240" -- 2DA6
           ,x"007f" -- 2DA8
           ,x"c800" -- 2DAA
           ,x"ed34" -- 2DAC
           ,x"75d7" -- 2DAE
           ,x"045b" -- 2DB0
           ,x"0420" -- 2DB2
           ,x"8d70" -- 2DB4
           ,x"0001" -- 2DB6
           ,x"0420" -- 2DB8
           ,x"b4e8" -- 2DBA
           ,x"10fa" -- 2DBC
           ,x"101e" -- 2DBE
           ,x"0420" -- 2DC0
           ,x"b526" -- 2DC2
           ,x"0280" -- 2DC4
           ,x"5600" -- 2DC6
           ,x"161c" -- 2DC8
           ,x"c0c2" -- 2DCA
           ,x"06a0" -- 2DCC
           ,x"b52a" -- 2DCE
           ,x"1007" -- 2DD0
           ,x"0420" -- 2DD2
           ,x"b540" -- 2DD4
           ,x"ccf2" -- 2DD6
           ,x"ccf2" -- 2DD8
           ,x"c4d2" -- 2DDA
           ,x"0460" -- 2DDC
           ,x"aefc" -- 2DDE
           ,x"0420" -- 2DE0
           ,x"b4e8" -- 2DE2
           ,x"1004" -- 2DE4
           ,x"1003" -- 2DE6
           ,x"0420" -- 2DE8
           ,x"8d70" -- 2DEA
           ,x"0001" -- 2DEC
           ,x"c102" -- 2DEE
           ,x"0280" -- 2DF0
           ,x"3f00" -- 2DF2
           ,x"1363" -- 2DF4
           ,x"0420" -- 2DF6
           ,x"8d70" -- 2DF8
           ,x"0007" -- 2DFA
           ,x"0280" -- 2DFC
           ,x"5600" -- 2DFE
           ,x"130e" -- 2E00
           ,x"0420" -- 2E02
           ,x"8d70" -- 2E04
           ,x"0024" -- 2E06
           ,x"c820" -- 2E08
           ,x"801a" -- 2E0A
           ,x"ef9e" -- 2E0C
           ,x"0420" -- 2E0E
           ,x"b558" -- 2E10
           ,x"06c1" -- 2E12
           ,x"ddc1" -- 2E14
           ,x"0280" -- 2E16
           ,x"4200" -- 2E18
           ,x"13f6" -- 2E1A
           ,x"10df" -- 2E1C
           ,x"c1c2" -- 2E1E
           ,x"0420" -- 2E20
           ,x"b4e8" -- 2E22
           ,x"1023" -- 2E24
           ,x"1022" -- 2E26
           ,x"d038" -- 2E28
           ,x"0280" -- 2E2A
           ,x"4200" -- 2E2C
           ,x"13ec" -- 2E2E
           ,x"0280" -- 2E30
           ,x"5e00" -- 2E32
           ,x"1357" -- 2E34
           ,x"0280" -- 2E36
           ,x"3e00" -- 2E38
           ,x"160d" -- 2E3A
           ,x"0420" -- 2E3C
           ,x"b4e8" -- 2E3E
           ,x"1004" -- 2E40
           ,x"1003" -- 2E42
           ,x"0420" -- 2E44
           ,x"8d70" -- 2E46
           ,x"000e" -- 2E48
           ,x"0280" -- 2E4A
           ,x"3f00" -- 2E4C
           ,x"16d3" -- 2E4E
           ,x"c802" -- 2E50
           ,x"ed3a" -- 2E52
           ,x"1001" -- 2E54
           ,x"0608" -- 2E56
           ,x"0420" -- 2E58
           ,x"b540" -- 2E5A
           ,x"c802" -- 2E5C
           ,x"ef9e" -- 2E5E
           ,x"0420" -- 2E60
           ,x"b05e" -- 2E62
           ,x"04e0" -- 2E64
           ,x"ed3a" -- 2E66
           ,x"75d7" -- 2E68
           ,x"10b8" -- 2E6A
           ,x"0705" -- 2E6C
           ,x"0280" -- 2E6E
           ,x"4000" -- 2E70
           ,x"1305" -- 2E72
           ,x"04c5" -- 2E74
           ,x"0280" -- 2E76
           ,x"3f00" -- 2E78
           ,x"1609" -- 2E7A
           ,x"0585" -- 2E7C
           ,x"c820" -- 2E7E
           ,x"801a" -- 2E80
           ,x"ef9e" -- 2E82
           ,x"0420" -- 2E84
           ,x"b558" -- 2E86
           ,x"c041" -- 2E88
           ,x"1505" -- 2E8A
           ,x"10a7" -- 2E8C
           ,x"c060" -- 2E8E
           ,x"ed04" -- 2E90
           ,x"6047" -- 2E92
           ,x"0601" -- 2E94
           ,x"c0c7" -- 2E96
           ,x"d132" -- 2E98
           ,x"1602" -- 2E9A
           ,x"c145" -- 2E9C
           ,x"1307" -- 2E9E
           ,x"ddc4" -- 2EA0
           ,x"81c2" -- 2EA2
           ,x"1402" -- 2EA4
           ,x"80c2" -- 2EA6
           ,x"1402" -- 2EA8
           ,x"0601" -- 2EAA
           ,x"16f5" -- 2EAC
           ,x"0915" -- 2EAE
           ,x"1601" -- 2EB0
           ,x"75d7" -- 2EB2
           ,x"0280" -- 2EB4
           ,x"5d00" -- 2EB6
           ,x"1639" -- 2EB8
           ,x"10b2" -- 2EBA
           ,x"0420" -- 2EBC
           ,x"b526" -- 2EBE
           ,x"04d2" -- 2EC0
           ,x"c1c4" -- 2EC2
           ,x"0420" -- 2EC4
           ,x"b288" -- 2EC6
           ,x"1007" -- 2EC8
           ,x"04c1" -- 2ECA
           ,x"1000" -- 2ECC
           ,x"d480" -- 2ECE
           ,x"04f3" -- 2ED0
           ,x"ccc1" -- 2ED2
           ,x"04d3" -- 2ED4
           ,x"102a" -- 2ED6
           ,x"d480" -- 2ED8
           ,x"c803" -- 2EDA
           ,x"ef7e" -- 2EDC
           ,x"0420" -- 2EDE
           ,x"bc32" -- 2EE0
           ,x"1024" -- 2EE2
           ,x"0420" -- 2EE4
           ,x"b4e8" -- 2EE6
           ,x"100e" -- 2EE8
           ,x"100d" -- 2EEA
           ,x"c820" -- 2EEC
           ,x"801a" -- 2EEE
           ,x"ef9e" -- 2EF0
           ,x"0420" -- 2EF2
           ,x"b558" -- 2EF4
           ,x"0601" -- 2EF6
           ,x"1103" -- 2EF8
           ,x"d032" -- 2EFA
           ,x"16fc" -- 2EFC
           ,x"0602" -- 2EFE
           ,x"ddf2" -- 2F00
           ,x"16fe" -- 2F02
           ,x"1013" -- 2F04
           ,x"c0c2" -- 2F06
           ,x"0701" -- 2F08
           ,x"0581" -- 2F0A
           ,x"d033" -- 2F0C
           ,x"16fd" -- 2F0E
           ,x"04c3" -- 2F10
           ,x"0583" -- 2F12
           ,x"d037" -- 2F14
           ,x"16fd" -- 2F16
           ,x"c107" -- 2F18
           ,x"a101" -- 2F1A
           ,x"0607" -- 2F1C
           ,x"0604" -- 2F1E
           ,x"d517" -- 2F20
           ,x"0603" -- 2F22
           ,x"15fb" -- 2F24
           ,x"ddf2" -- 2F26
           ,x"0601" -- 2F28
           ,x"15fd" -- 2F2A
           ,x"0460" -- 2F2C
           ,x"aefc" -- 2F2E
           ,x"c28b" -- 2F30
           ,x"0420" -- 2F32
           ,x"be74" -- 2F34
           ,x"c101" -- 2F36
           ,x"06a0" -- 2F38
           ,x"bbd6" -- 2F3A
           ,x"c084" -- 2F3C
           ,x"c101" -- 2F3E
           ,x"06a0" -- 2F40
           ,x"bbd6" -- 2F42
           ,x"c081" -- 2F44
           ,x"c07a" -- 2F46
           ,x"0203" -- 2F48
           ,x"045a" -- 2F4A
           ,x"0441" -- 2F4C
           ,x"06a0" -- 2F4E
           ,x"9930" -- 2F50
           ,x"0264" -- 2F52
           ,x"1008" -- 2F54
           ,x"06a0" -- 2F56
           ,x"9930" -- 2F58
           ,x"045a" -- 2F5A
           ,x"2902" -- 2F5C
           ,x"1003" -- 2F5E
           ,x"06a0" -- 2F60
           ,x"9930" -- 2F62
           ,x"0244" -- 2F64
           ,x"c804" -- 2F66
           ,x"ef6a" -- 2F68
           ,x"0202" -- 2F6A
           ,x"ef68" -- 2F6C
           ,x"0460" -- 2F6E
           ,x"b82e" -- 2F70
           ,x"0420" -- 2F72
           ,x"be74" -- 2F74
           ,x"c081" -- 2F76
           ,x"06a0" -- 2F78
           ,x"bbd6" -- 2F7A
           ,x"0541" -- 2F7C
           ,x"c801" -- 2F7E
           ,x"ef6a" -- 2F80
           ,x"10f3" -- 2F82
           ,x"9838" -- 2F84
           ,x"ad1f" -- 2F86
           ,x"160a" -- 2F88
           ,x"0420" -- 2F8A
           ,x"b540" -- 2F8C
           ,x"06a0" -- 2F8E
           ,x"bc16" -- 2F90
           ,x"06a0" -- 2F92
           ,x"c1ba" -- 2F94
           ,x"06c3" -- 2F96
           ,x"d443" -- 2F98
           ,x"0460" -- 2F9A
           ,x"aefc" -- 2F9C
           ,x"0460" -- 2F9E
           ,x"97b2" -- 2FA0
           ,x"06a0" -- 2FA2
           ,x"bc16" -- 2FA4
           ,x"d051" -- 2FA6
           ,x"0981" -- 2FA8
           ,x"0420" -- 2FAA
           ,x"be74" -- 2FAC
           ,x"c801" -- 2FAE
           ,x"ef6a" -- 2FB0
           ,x"0460" -- 2FB2
           ,x"b6be" -- 2FB4
           ,x"d052" -- 2FB6
           ,x"10f7" -- 2FB8
           ,x"04c3" -- 2FBA
           ,x"d5f2" -- 2FBC
           ,x"130d" -- 2FBE
           ,x"9817" -- 2FC0
           ,x"c84f" -- 2FC2
           ,x"130b" -- 2FC4
           ,x"0587" -- 2FC6
           ,x"c2a0" -- 2FC8
           ,x"ed04" -- 2FCA
           ,x"060a" -- 2FCC
           ,x"8287" -- 2FCE
           ,x"1303" -- 2FD0
           ,x"0605" -- 2FD2
           ,x"15f3" -- 2FD4
           ,x"05cb" -- 2FD6
           ,x"75d7" -- 2FD8
           ,x"045b" -- 2FDA
           ,x"04c1" -- 2FDC
           ,x"c282" -- 2FDE
           ,x"04c0" -- 2FE0
           ,x"d03a" -- 2FE2
           ,x"0220" -- 2FE4
           ,x"d000" -- 2FE6
           ,x"110e" -- 2FE8
           ,x"0280" -- 2FEA
           ,x"0900" -- 2FEC
           ,x"1208" -- 2FEE
           ,x"0220" -- 2FF0
           ,x"f900" -- 2FF2
           ,x"0280" -- 2FF4
           ,x"0a00" -- 2FF6
           ,x"1106" -- 2FF8
           ,x"0280" -- 2FFA
           ,x"0f00" -- 2FFC
           ,x"1b03" -- 2FFE
           ,x"0a41" -- 3000
           ,x"b040" -- 3002
           ,x"10ed" -- 3004
           ,x"0280" -- 3006
           ,x"0700" -- 3008
           ,x"16dd" -- 300A
           ,x"d041" -- 300C
           ,x"13db" -- 300E
           ,x"c08a" -- 3010
           ,x"d5c1" -- 3012
           ,x"9801" -- 3014
           ,x"c0ea" -- 3016
           ,x"16d6" -- 3018
           ,x"0643" -- 301A
           ,x"10d4" -- 301C
           ,x"9838" -- 301E
           ,x"ad1f" -- 3020
           ,x"1609" -- 3022
           ,x"0420" -- 3024
           ,x"b540" -- 3026
           ,x"06a0" -- 3028
           ,x"bc16" -- 302A
           ,x"06a0" -- 302C
           ,x"c1ba" -- 302E
           ,x"c443" -- 3030
           ,x"0460" -- 3032
           ,x"aefc" -- 3034
           ,x"0460" -- 3036
           ,x"97b2" -- 3038
           ,x"06a0" -- 303A
           ,x"bc16" -- 303C
           ,x"c051" -- 303E
           ,x"0420" -- 3040
           ,x"be74" -- 3042
           ,x"c801" -- 3044
           ,x"ef6a" -- 3046
           ,x"0460" -- 3048
           ,x"b6be" -- 304A
           ,x"c042" -- 304C
           ,x"10fa" -- 304E
           ,x"06a0" -- 3050
           ,x"a364" -- 3052
           ,x"d018" -- 3054
           ,x"1313" -- 3056
           ,x"c820" -- 3058
           ,x"8008" -- 305A
           ,x"ef9e" -- 305C
           ,x"0420" -- 305E
           ,x"b558" -- 3060
           ,x"0280" -- 3062
           ,x"3f00" -- 3064
           ,x"160f" -- 3066
           ,x"c820" -- 3068
           ,x"801a" -- 306A
           ,x"ef9e" -- 306C
           ,x"0420" -- 306E
           ,x"b558" -- 3070
           ,x"c801" -- 3072
           ,x"ede0" -- 3074
           ,x"6801" -- 3076
           ,x"edee" -- 3078
           ,x"0460" -- 307A
           ,x"8124" -- 307C
           ,x"0201" -- 307E
           ,x"0064" -- 3080
           ,x"c801" -- 3082
           ,x"edee" -- 3084
           ,x"0201" -- 3086
           ,x"000a" -- 3088
           ,x"10f3" -- 308A
           ,x"c820" -- 308C
           ,x"801a" -- 308E
           ,x"ef9e" -- 3090
           ,x"0420" -- 3092
           ,x"b558" -- 3094
           ,x"0280" -- 3096
           ,x"3b00" -- 3098
           ,x"1614" -- 309A
           ,x"04c2" -- 309C
           ,x"d0b8" -- 309E
           ,x"0972" -- 30A0
           ,x"c0c2" -- 30A2
           ,x"0643" -- 30A4
           ,x"1303" -- 30A6
           ,x"0223" -- 30A8
           ,x"fffd" -- 30AA
           ,x"150b" -- 30AC
           ,x"0601" -- 30AE
           ,x"1105" -- 30B0
           ,x"1306" -- 30B2
           ,x"05c8" -- 30B4
           ,x"9838" -- 30B6
           ,x"c8c0" -- 30B8
           ,x"13f9" -- 30BA
           ,x"0460" -- 30BC
           ,x"af02" -- 30BE
           ,x"0460" -- 30C0
           ,x"952a" -- 30C2
           ,x"0460" -- 30C4
           ,x"97b2" -- 30C6
           ,x"0420" -- 30C8
           ,x"b4e8" -- 30CA
           ,x"1032" -- 30CC
           ,x"1031" -- 30CE
           ,x"9838" -- 30D0
           ,x"baa2" -- 30D2
           ,x"1649" -- 30D4
           ,x"c820" -- 30D6
           ,x"801e" -- 30D8
           ,x"ef9e" -- 30DA
           ,x"0420" -- 30DC
           ,x"b558" -- 30DE
           ,x"c820" -- 30E0
           ,x"801a" -- 30E2
           ,x"ef9e" -- 30E4
           ,x"0420" -- 30E6
           ,x"b558" -- 30E8
           ,x"0280" -- 30EA
           ,x"4d00" -- 30EC
           ,x"163c" -- 30EE
           ,x"0281" -- 30F0
           ,x"0017" -- 30F2
           ,x"1b39" -- 30F4
           ,x"0283" -- 30F6
           ,x"0027" -- 30F8
           ,x"1b36" -- 30FA
           ,x"c2a0" -- 30FC
           ,x"804c" -- 30FE
           ,x"1305" -- 3100
           ,x"0283" -- 3102
           ,x"001f" -- 3104
           ,x"1b30" -- 3106
           ,x"0a31" -- 3108
           ,x"0a33" -- 310A
           ,x"06c1" -- 310C
           ,x"06c3" -- 310E
           ,x"c020" -- 3110
           ,x"ed36" -- 3112
           ,x"1603" -- 3114
           ,x"0420" -- 3116
           ,x"818c" -- 3118
           ,x"1d00" -- 311A
           ,x"d803" -- 311C
           ,x"ef42" -- 311E
           ,x"d801" -- 3120
           ,x"ef43" -- 3122
           ,x"c800" -- 3124
           ,x"ed36" -- 3126
           ,x"162b" -- 3128
           ,x"0420" -- 312A
           ,x"818c" -- 312C
           ,x"1c00" -- 312E
           ,x"1027" -- 3130
           ,x"c0c7" -- 3132
           ,x"c1c2" -- 3134
           ,x"0201" -- 3136
           ,x"0001" -- 3138
           ,x"0420" -- 313A
           ,x"b284" -- 313C
           ,x"1014" -- 313E
           ,x"0587" -- 3140
           ,x"c141" -- 3142
           ,x"d000" -- 3144
           ,x"130d" -- 3146
           ,x"0202" -- 3148
           ,x"9cb4" -- 314A
           ,x"c132" -- 314C
           ,x"130c" -- 314E
           ,x"9100" -- 3150
           ,x"16fc" -- 3152
           ,x"06c4" -- 3154
           ,x"d004" -- 3156
           ,x"0420" -- 3158
           ,x"816c" -- 315A
           ,x"0605" -- 315C
           ,x"16fb" -- 315E
           ,x"10ea" -- 3160
           ,x"0608" -- 3162
           ,x"c1c3" -- 3164
           ,x"100c" -- 3166
           ,x"0420" -- 3168
           ,x"8d70" -- 316A
           ,x"000f" -- 316C
           ,x"020e" -- 316E
           ,x"0084" -- 3170
           ,x"c020" -- 3172
           ,x"ede4" -- 3174
           ,x"1601" -- 3176
           ,x"093e" -- 3178
           ,x"c1e0" -- 317A
           ,x"ed04" -- 317C
           ,x"070f" -- 317E
           ,x"058f" -- 3180
           ,x"06a0" -- 3182
           ,x"8724" -- 3184
           ,x"1b00" -- 3186
           ,x"1b3c" -- 3188
           ,x"1b47" -- 318A
           ,x"1d3e" -- 318C
           ,x"583f" -- 318E
           ,x"6040" -- 3190
           ,x"6739" -- 3192
           ,x"a13d" -- 3194
           ,x"0000" -- 3196
           ,x"0608" -- 3198
           ,x"0420" -- 319A
           ,x"b4e8" -- 319C
           ,x"103c" -- 319E
           ,x"103b" -- 31A0
           ,x"0420" -- 31A2
           ,x"b540" -- 31A4
           ,x"c120" -- 31A6
           ,x"ed3a" -- 31A8
           ,x"1602" -- 31AA
           ,x"dde0" -- 31AC
           ,x"c0e4" -- 31AE
           ,x"c802" -- 31B0
           ,x"ef9e" -- 31B2
           ,x"0420" -- 31B4
           ,x"b05e" -- 31B6
           ,x"0608" -- 31B8
           ,x"10e1" -- 31BA
           ,x"0460" -- 31BC
           ,x"977e" -- 31BE
           ,x"0420" -- 31C0
           ,x"b4e8" -- 31C2
           ,x"1026" -- 31C4
           ,x"1025" -- 31C6
           ,x"0202" -- 31C8
           ,x"0005" -- 31CA
           ,x"9818" -- 31CC
           ,x"c8c0" -- 31CE
           ,x"1607" -- 31D0
           ,x"0588" -- 31D2
           ,x"c820" -- 31D4
           ,x"801a" -- 31D6
           ,x"ef9e" -- 31D8
           ,x"0420" -- 31DA
           ,x"b558" -- 31DC
           ,x"100b" -- 31DE
           ,x"9818" -- 31E0
           ,x"c8e0" -- 31E2
           ,x"160c" -- 31E4
           ,x"0588" -- 31E6
           ,x"c820" -- 31E8
           ,x"801a" -- 31EA
           ,x"ef9e" -- 31EC
           ,x"0420" -- 31EE
           ,x"b558" -- 31F0
           ,x"0642" -- 31F2
           ,x"0a81" -- 31F4
           ,x"06a0" -- 31F6
           ,x"9ca8" -- 31F8
           ,x"0607" -- 31FA
           ,x"10dd" -- 31FC
           ,x"c820" -- 31FE
           ,x"801a" -- 3200
           ,x"ef9e" -- 3202
           ,x"0420" -- 3204
           ,x"b558" -- 3206
           ,x"dde0" -- 3208
           ,x"c0e4" -- 320A
           ,x"06a0" -- 320C
           ,x"9c8e" -- 320E
           ,x"10d3" -- 3210
           ,x"c802" -- 3212
           ,x"ed3a" -- 3214
           ,x"10d0" -- 3216
           ,x"c14e" -- 3218
           ,x"a160" -- 321A
           ,x"ed04" -- 321C
           ,x"6147" -- 321E
           ,x"06a0" -- 3220
           ,x"99ba" -- 3222
           ,x"1005" -- 3224
           ,x"06a0" -- 3226
           ,x"9772" -- 3228
           ,x"a803" -- 322A
           ,x"ed34" -- 322C
           ,x"10f4" -- 322E
           ,x"a803" -- 3230
           ,x"ed34" -- 3232
           ,x"10c1" -- 3234
           ,x"06a0" -- 3236
           ,x"9c82" -- 3238
           ,x"0240" -- 323A
           ,x"0007" -- 323C
           ,x"0220" -- 323E
           ,x"fff8" -- 3240
           ,x"06a0" -- 3242
           ,x"9c78" -- 3244
           ,x"06a0" -- 3246
           ,x"9c82" -- 3248
           ,x"600e" -- 324A
           ,x"1199" -- 324C
           ,x"06a0" -- 324E
           ,x"9772" -- 3250
           ,x"1096" -- 3252
           ,x"c820" -- 3254
           ,x"801a" -- 3256
           ,x"ef9e" -- 3258
           ,x"0420" -- 325A
           ,x"b558" -- 325C
           ,x"0608" -- 325E
           ,x"0241" -- 3260
           ,x"007f" -- 3262
           ,x"06a0" -- 3264
           ,x"9c82" -- 3266
           ,x"6001" -- 3268
           ,x"158a" -- 326A
           ,x"c060" -- 326C
           ,x"ede4" -- 326E
           ,x"1387" -- 3270
           ,x"06a0" -- 3272
           ,x"9c78" -- 3274
           ,x"1084" -- 3276
           ,x"0580" -- 3278
           ,x"1508" -- 327A
           ,x"dde0" -- 327C
           ,x"c0e4" -- 327E
           ,x"10fb" -- 3280
           ,x"c020" -- 3282
           ,x"ed34" -- 3284
           ,x"a007" -- 3286
           ,x"6020" -- 3288
           ,x"ed04" -- 328A
           ,x"045b" -- 328C
           ,x"04c0" -- 328E
           ,x"dde0" -- 3290
           ,x"9cc4" -- 3292
           ,x"0202" -- 3294
           ,x"0004" -- 3296
           ,x"c101" -- 3298
           ,x"0a41" -- 329A
           ,x"09c4" -- 329C
           ,x"1602" -- 329E
           ,x"c000" -- 32A0
           ,x"1303" -- 32A2
           ,x"dde4" -- 32A4
           ,x"9cc4" -- 32A6
           ,x"0700" -- 32A8
           ,x"0602" -- 32AA
           ,x"15f5" -- 32AC
           ,x"dde0" -- 32AE
           ,x"9cc0" -- 32B0
           ,x"045b" -- 32B2
           ,x"550b" -- 32B4
           ,x"440a" -- 32B6
           ,x"4c08" -- 32B8
           ,x"5209" -- 32BA
           ,x"420d" -- 32BC
           ,x"430c" -- 32BE
           ,x"481e" -- 32C0
           ,x"0000" -- 32C2
           ,x"3031" -- 32C4
           ,x"3233" -- 32C6
           ,x"3435" -- 32C8
           ,x"3637" -- 32CA
           ,x"3839" -- 32CC
           ,x"4142" -- 32CE
           ,x"4344" -- 32D0
           ,x"4546" -- 32D2
           ,x"06a0" -- 32D4
           ,x"a364" -- 32D6
           ,x"c0a0" -- 32D8
           ,x"ede6" -- 32DA
           ,x"1303" -- 32DC
           ,x"c822" -- 32DE
           ,x"fffa" -- 32E0
           ,x"ed32" -- 32E2
           ,x"c820" -- 32E4
           ,x"801a" -- 32E6
           ,x"ef9e" -- 32E8
           ,x"0420" -- 32EA
           ,x"b558" -- 32EC
           ,x"0280" -- 32EE
           ,x"3800" -- 32F0
           ,x"1621" -- 32F2
           ,x"c820" -- 32F4
           ,x"801e" -- 32F6
           ,x"ef9e" -- 32F8
           ,x"0420" -- 32FA
           ,x"b558" -- 32FC
           ,x"c3c3" -- 32FE
           ,x"c3a0" -- 3300
           ,x"edd4" -- 3302
           ,x"064e" -- 3304
           ,x"880e" -- 3306
           ,x"edd2" -- 3308
           ,x"1213" -- 330A
           ,x"022e" -- 330C
           ,x"fffc" -- 330E
           ,x"8781" -- 3310
           ,x"15f9" -- 3312
           ,x"880e" -- 3314
           ,x"edd2" -- 3316
           ,x"1a0c" -- 3318
           ,x"83de" -- 331A
           ,x"150a" -- 331C
           ,x"04c0" -- 331E
           ,x"c05e" -- 3320
           ,x"0720" -- 3322
           ,x"8046" -- 3324
           ,x"06a0" -- 3326
           ,x"a77c" -- 3328
           ,x"0420" -- 332A
           ,x"8194" -- 332C
           ,x"10e8" -- 332E
           ,x"10e7" -- 3330
           ,x"0460" -- 3332
           ,x"8116" -- 3334
           ,x"0460" -- 3336
           ,x"aef2" -- 3338
           ,x"0240" -- 333A
           ,x"ff00" -- 333C
           ,x"0280" -- 333E
           ,x"0d00" -- 3340
           ,x"1602" -- 3342
           ,x"75d7" -- 3344
           ,x"045b" -- 3346
           ,x"0280" -- 3348
           ,x"2000" -- 334A
           ,x"1402" -- 334C
           ,x"046b" -- 334E
           ,x"0002" -- 3350
           ,x"0280" -- 3352
           ,x"7f00" -- 3354
           ,x"1605" -- 3356
           ,x"0584" -- 3358
           ,x"8807" -- 335A
           ,x"ed04" -- 335C
           ,x"1b06" -- 335E
           ,x"1011" -- 3360
           ,x"8807" -- 3362
           ,x"ed0c" -- 3364
           ,x"14fc" -- 3366
           ,x"ddc0" -- 3368
           ,x"100c" -- 336A
           ,x"0607" -- 336C
           ,x"0584" -- 336E
           ,x"0620" -- 3370
           ,x"ed34" -- 3372
           ,x"0420" -- 3374
           ,x"818c" -- 3376
           ,x"0800" -- 3378
           ,x"0420" -- 337A
           ,x"818c" -- 337C
           ,x"2000" -- 337E
           ,x"0200" -- 3380
           ,x"0800" -- 3382
           ,x"046b" -- 3384
           ,x"0004" -- 3386
           ,x"c820" -- 3388
           ,x"8006" -- 338A
           ,x"ef9e" -- 338C
           ,x"0420" -- 338E
           ,x"b558" -- 3390
           ,x"0460" -- 3392
           ,x"aefc" -- 3394
           ,x"c188" -- 3396
           ,x"c160" -- 3398
           ,x"ede8" -- 339A
           ,x"c220" -- 339C
           ,x"edec" -- 339E
           ,x"1309" -- 33A0
           ,x"04c0" -- 33A2
           ,x"d038" -- 33A4
           ,x"1306" -- 33A6
           ,x"0280" -- 33A8
           ,x"3f00" -- 33AA
           ,x"1312" -- 33AC
           ,x"0420" -- 33AE
           ,x"8d70" -- 33B0
           ,x"0017" -- 33B2
           ,x"c220" -- 33B4
           ,x"edea" -- 33B6
           ,x"0228" -- 33B8
           ,x"fffc" -- 33BA
           ,x"8808" -- 33BC
           ,x"edd2" -- 33BE
           ,x"1af6" -- 33C0
           ,x"c808" -- 33C2
           ,x"edea" -- 33C4
           ,x"c218" -- 33C6
           ,x"a220" -- 33C8
           ,x"ed0e" -- 33CA
           ,x"9838" -- 33CC
           ,x"b052" -- 33CE
           ,x"16f1" -- 33D0
           ,x"0420" -- 33D2
           ,x"b4e8" -- 33D4
           ,x"1004" -- 33D6
           ,x"1003" -- 33D8
           ,x"0420" -- 33DA
           ,x"b540" -- 33DC
           ,x"05cb" -- 33DE
           ,x"0608" -- 33E0
           ,x"c808" -- 33E2
           ,x"edec" -- 33E4
           ,x"c206" -- 33E6
           ,x"c805" -- 33E8
           ,x"ede8" -- 33EA
           ,x"045b" -- 33EC
           ,x"0420" -- 33EE
           ,x"8d70" -- 33F0
           ,x"0018" -- 33F2
           ,x"0420" -- 33F4
           ,x"b4e8" -- 33F6
           ,x"10fa" -- 33F8
           ,x"1010" -- 33FA
           ,x"0420" -- 33FC
           ,x"b526" -- 33FE
           ,x"c1c2" -- 3400
           ,x"06a0" -- 3402
           ,x"9d96" -- 3404
           ,x"10f3" -- 3406
           ,x"cdf2" -- 3408
           ,x"cdf2" -- 340A
           ,x"c5d2" -- 340C
           ,x"c020" -- 340E
           ,x"ede8" -- 3410
           ,x"0280" -- 3412
           ,x"3f00" -- 3414
           ,x"13ee" -- 3416
           ,x"0460" -- 3418
           ,x"aefc" -- 341A
           ,x"c1c2" -- 341C
           ,x"06a0" -- 341E
           ,x"9d96" -- 3420
           ,x"1001" -- 3422
           ,x"10e4" -- 3424
           ,x"0205" -- 3426
           ,x"0084" -- 3428
           ,x"06a0" -- 342A
           ,x"99ba" -- 342C
           ,x"10ef" -- 342E
           ,x"06a0" -- 3430
           ,x"aeb2" -- 3432
           ,x"06a0" -- 3434
           ,x"b52a" -- 3436
           ,x"100e" -- 3438
           ,x"c820" -- 343A
           ,x"801a" -- 343C
           ,x"ef9e" -- 343E
           ,x"0420" -- 3440
           ,x"b558" -- 3442
           ,x"c088" -- 3444
           ,x"06a0" -- 3446
           ,x"a2a6" -- 3448
           ,x"8e38" -- 344A
           ,x"c808" -- 344C
           ,x"edea" -- 344E
           ,x"c202" -- 3450
           ,x"0460" -- 3452
           ,x"aefc" -- 3454
           ,x"0460" -- 3456
           ,x"aef8" -- 3458
           ,x"0001" -- 345A
           ,x"0002" -- 345C
           ,x"000f" -- 345E
           ,x"0040" -- 3460
           ,x"000d" -- 3462
           ,x"0009" -- 3464
           ,x"0004" -- 3466
           ,x"0041" -- 3468
           ,x"0003" -- 346A
           ,x"4544" -- 346C
           ,x"476d" -- 346E
           ,x"6e6f" -- 3470
           ,x"3c3e" -- 3472
           ,x"3f41" -- 3474
           ,x"403a" -- 3476
           ,x"3b00" -- 3478
           ,x"06a0" -- 347A
           ,x"a364" -- 347C
           ,x"0201" -- 347E
           ,x"000a" -- 3480
           ,x"c081" -- 3482
           ,x"9838" -- 3484
           ,x"9e77" -- 3486
           ,x"130c" -- 3488
           ,x"0608" -- 348A
           ,x"06a0" -- 348C
           ,x"b52a" -- 348E
           ,x"100d" -- 3490
           ,x"c820" -- 3492
           ,x"801c" -- 3494
           ,x"ef9e" -- 3496
           ,x"0420" -- 3498
           ,x"b558" -- 349A
           ,x"9800" -- 349C
           ,x"9e77" -- 349E
           ,x"1605" -- 34A0
           ,x"c820" -- 34A2
           ,x"801a" -- 34A4
           ,x"ef9e" -- 34A6
           ,x"0420" -- 34A8
           ,x"b558" -- 34AA
           ,x"c801" -- 34AC
           ,x"ed1c" -- 34AE
           ,x"6081" -- 34B0
           ,x"c802" -- 34B2
           ,x"ed1a" -- 34B4
           ,x"0720" -- 34B6
           ,x"8046" -- 34B8
           ,x"06a0" -- 34BA
           ,x"a128" -- 34BC
           ,x"0000" -- 34BE
           ,x"c120" -- 34C0
           ,x"edd8" -- 34C2
           ,x"c1a0" -- 34C4
           ,x"edda" -- 34C6
           ,x"0226" -- 34C8
           ,x"fffa" -- 34CA
           ,x"c0a0" -- 34CC
           ,x"ed1a" -- 34CE
           ,x"c160" -- 34D0
           ,x"edd4" -- 34D2
           ,x"0645" -- 34D4
           ,x"0645" -- 34D6
           ,x"8160" -- 34D8
           ,x"edd2" -- 34DA
           ,x"1a57" -- 34DC
           ,x"04d4" -- 34DE
           ,x"c1e0" -- 34E0
           ,x"ed1a" -- 34E2
           ,x"c160" -- 34E4
           ,x"edd4" -- 34E6
           ,x"0645" -- 34E8
           ,x"a1e0" -- 34EA
           ,x"ed1c" -- 34EC
           ,x"0225" -- 34EE
           ,x"fffc" -- 34F0
           ,x"8805" -- 34F2
           ,x"edd2" -- 34F4
           ,x"1a11" -- 34F6
           ,x"c120" -- 34F8
           ,x"edd8" -- 34FA
           ,x"c514" -- 34FC
           ,x"130b" -- 34FE
           ,x"8d15" -- 3500
           ,x"1607" -- 3502
           ,x"0644" -- 3504
           ,x"0534" -- 3506
           ,x"c014" -- 3508
           ,x"dc07" -- 350A
           ,x"06c7" -- 350C
           ,x"d407" -- 350E
           ,x"06c7" -- 3510
           ,x"05c4" -- 3512
           ,x"10f3" -- 3514
           ,x"c547" -- 3516
           ,x"10e8" -- 3518
           ,x"c120" -- 351A
           ,x"edd8" -- 351C
           ,x"c014" -- 351E
           ,x"112d" -- 3520
           ,x"132f" -- 3522
           ,x"c064" -- 3524
           ,x"0002" -- 3526
           ,x"c160" -- 3528
           ,x"edd2" -- 352A
           ,x"c0b5" -- 352C
           ,x"c235" -- 352E
           ,x"a220" -- 3530
           ,x"ed0e" -- 3532
           ,x"8201" -- 3534
           ,x"1afa" -- 3536
           ,x"06a0" -- 3538
           ,x"a226" -- 353A
           ,x"0d0a" -- 353C
           ,x"4261" -- 353E
           ,x"6420" -- 3540
           ,x"6c69" -- 3542
           ,x"6e65" -- 3544
           ,x"206e" -- 3546
           ,x"6f2e" -- 3548
           ,x"20d8" -- 354A
           ,x"c820" -- 354C
           ,x"8018" -- 354E
           ,x"ef9e" -- 3550
           ,x"0420" -- 3552
           ,x"b05a" -- 3554
           ,x"06a0" -- 3556
           ,x"a22a" -- 3558
           ,x"2920" -- 355A
           ,x"696e" -- 355C
           ,x"206e" -- 355E
           ,x"6577" -- 3560
           ,x"206c" -- 3562
           ,x"696e" -- 3564
           ,x"65e0" -- 3566
           ,x"c820" -- 3568
           ,x"801c" -- 356A
           ,x"ef9e" -- 356C
           ,x"0420" -- 356E
           ,x"b05a" -- 3570
           ,x"06a0" -- 3572
           ,x"a22a" -- 3574
           ,x"0000" -- 3576
           ,x"0420" -- 3578
           ,x"8174" -- 357A
           ,x"04f4" -- 357C
           ,x"04f4" -- 357E
           ,x"10ce" -- 3580
           ,x"06a0" -- 3582
           ,x"a128" -- 3584
           ,x"0009" -- 3586
           ,x"0460" -- 3588
           ,x"8124" -- 358A
           ,x"a0a0" -- 358C
           ,x"ed1c" -- 358E
           ,x"c215" -- 3590
           ,x"a220" -- 3592
           ,x"ed0e" -- 3594
           ,x"d618" -- 3596
           ,x"139d" -- 3598
           ,x"d0d8" -- 359A
           ,x"9818" -- 359C
           ,x"9e5b" -- 359E
           ,x"1308" -- 35A0
           ,x"9818" -- 35A2
           ,x"9e5d" -- 35A4
           ,x"1305" -- 35A6
           ,x"1012" -- 35A8
           ,x"0588" -- 35AA
           ,x"9818" -- 35AC
           ,x"9e6f" -- 35AE
           ,x"166e" -- 35B0
           ,x"0588" -- 35B2
           ,x"05c8" -- 35B4
           ,x"d618" -- 35B6
           ,x"1306" -- 35B8
           ,x"9818" -- 35BA
           ,x"9e72" -- 35BC
           ,x"1303" -- 35BE
           ,x"9818" -- 35C0
           ,x"9e6e" -- 35C2
           ,x"1664" -- 35C4
           ,x"0648" -- 35C6
           ,x"06a0" -- 35C8
           ,x"a108" -- 35CA
           ,x"1052" -- 35CC
           ,x"9818" -- 35CE
           ,x"9e5f" -- 35D0
           ,x"160d" -- 35D2
           ,x"0588" -- 35D4
           ,x"d618" -- 35D6
           ,x"134c" -- 35D8
           ,x"9818" -- 35DA
           ,x"9e72" -- 35DC
           ,x"1349" -- 35DE
           ,x"9818" -- 35E0
           ,x"9e6e" -- 35E2
           ,x"1346" -- 35E4
           ,x"9818" -- 35E6
           ,x"9e73" -- 35E8
           ,x"1343" -- 35EA
           ,x"10df" -- 35EC
           ,x"9818" -- 35EE
           ,x"9e61" -- 35F0
           ,x"1303" -- 35F2
           ,x"9818" -- 35F4
           ,x"9e69" -- 35F6
           ,x"1629" -- 35F8
           ,x"0588" -- 35FA
           ,x"9818" -- 35FC
           ,x"9e78" -- 35FE
           ,x"131a" -- 3600
           ,x"9818" -- 3602
           ,x"9e72" -- 3604
           ,x"1317" -- 3606
           ,x"9818" -- 3608
           ,x"9e6f" -- 360A
           ,x"1309" -- 360C
           ,x"9818" -- 360E
           ,x"9e70" -- 3610
           ,x"1306" -- 3612
           ,x"9818" -- 3614
           ,x"9e71" -- 3616
           ,x"1605" -- 3618
           ,x"0228" -- 361A
           ,x"0006" -- 361C
           ,x"10ed" -- 361E
           ,x"05c8" -- 3620
           ,x"10eb" -- 3622
           ,x"9818" -- 3624
           ,x"9e6c" -- 3626
           ,x"1303" -- 3628
           ,x"9818" -- 362A
           ,x"9e6d" -- 362C
           ,x"16e5" -- 362E
           ,x"d038" -- 3630
           ,x"16fe" -- 3632
           ,x"10e3" -- 3634
           ,x"0588" -- 3636
           ,x"9803" -- 3638
           ,x"9e69" -- 363A
           ,x"13ac" -- 363C
           ,x"0588" -- 363E
           ,x"06a0" -- 3640
           ,x"a108" -- 3642
           ,x"9818" -- 3644
           ,x"9e74" -- 3646
           ,x"1614" -- 3648
           ,x"10f9" -- 364A
           ,x"9818" -- 364C
           ,x"9e63" -- 364E
           ,x"130f" -- 3650
           ,x"9818" -- 3652
           ,x"9e65" -- 3654
           ,x"13a9" -- 3656
           ,x"9818" -- 3658
           ,x"9e67" -- 365A
           ,x"1603" -- 365C
           ,x"d038" -- 365E
           ,x"16fe" -- 3660
           ,x"1006" -- 3662
           ,x"9818" -- 3664
           ,x"9e6b" -- 3666
           ,x"1604" -- 3668
           ,x"0588" -- 366A
           ,x"1094" -- 366C
           ,x"05c8" -- 366E
           ,x"0588" -- 3670
           ,x"d618" -- 3672
           ,x"13fb" -- 3674
           ,x"9818" -- 3676
           ,x"9e72" -- 3678
           ,x"13f7" -- 367A
           ,x"9818" -- 367C
           ,x"9e75" -- 367E
           ,x"1618" -- 3680
           ,x"9803" -- 3682
           ,x"9e63" -- 3684
           ,x"1615" -- 3686
           ,x"0588" -- 3688
           ,x"9818" -- 368A
           ,x"9e6f" -- 368C
           ,x"1626" -- 368E
           ,x"0588" -- 3690
           ,x"05c8" -- 3692
           ,x"d618" -- 3694
           ,x"1397" -- 3696
           ,x"9818" -- 3698
           ,x"9e72" -- 369A
           ,x"1394" -- 369C
           ,x"9818" -- 369E
           ,x"9e6e" -- 36A0
           ,x"1391" -- 36A2
           ,x"9818" -- 36A4
           ,x"9e74" -- 36A6
           ,x"138e" -- 36A8
           ,x"9818" -- 36AA
           ,x"9e76" -- 36AC
           ,x"1616" -- 36AE
           ,x"108a" -- 36B0
           ,x"9818" -- 36B2
           ,x"9e6c" -- 36B4
           ,x"13d3" -- 36B6
           ,x"9818" -- 36B8
           ,x"9e6d" -- 36BA
           ,x"13d0" -- 36BC
           ,x"9818" -- 36BE
           ,x"9e6e" -- 36C0
           ,x"13cd" -- 36C2
           ,x"9818" -- 36C4
           ,x"9e6f" -- 36C6
           ,x"13d2" -- 36C8
           ,x"9818" -- 36CA
           ,x"9e70" -- 36CC
           ,x"13cf" -- 36CE
           ,x"9818" -- 36D0
           ,x"9e71" -- 36D2
           ,x"16cd" -- 36D4
           ,x"0228" -- 36D6
           ,x"0006" -- 36D8
           ,x"10cb" -- 36DA
           ,x"06a0" -- 36DC
           ,x"a226" -- 36DE
           ,x"0d0a" -- 36E0
           ,x"5072" -- 36E2
           ,x"6f62" -- 36E4
           ,x"6c65" -- 36E6
           ,x"6d20" -- 36E8
           ,x"7769" -- 36EA
           ,x"7468" -- 36EC
           ,x"206e" -- 36EE
           ,x"6577" -- 36F0
           ,x"206c" -- 36F2
           ,x"696e" -- 36F4
           ,x"65e0" -- 36F6
           ,x"c820" -- 36F8
           ,x"801c" -- 36FA
           ,x"ef9e" -- 36FC
           ,x"0420" -- 36FE
           ,x"b05a" -- 3700
           ,x"0420" -- 3702
           ,x"8174" -- 3704
           ,x"10b5" -- 3706
           ,x"8106" -- 3708
           ,x"1a06" -- 370A
           ,x"dd38" -- 370C
           ,x"dd18" -- 370E
           ,x"0608" -- 3710
           ,x"cd08" -- 3712
           ,x"05c8" -- 3714
           ,x"045b" -- 3716
           ,x"c120" -- 3718
           ,x"edd8" -- 371A
           ,x"05c6" -- 371C
           ,x"04f4" -- 371E
           ,x"8106" -- 3720
           ,x"14fd" -- 3722
           ,x"0460" -- 3724
           ,x"a5a6" -- 3726
           ,x"c83b" -- 3728
           ,x"ed14" -- 372A
           ,x"c80b" -- 372C
           ,x"ed16" -- 372E
           ,x"04e0" -- 3730
           ,x"ed18" -- 3732
           ,x"0720" -- 3734
           ,x"ede2" -- 3736
           ,x"c220" -- 3738
           ,x"edd4" -- 373A
           ,x"0648" -- 373C
           ,x"8808" -- 373E
           ,x"edd2" -- 3740
           ,x"120f" -- 3742
           ,x"0228" -- 3744
           ,x"fffc" -- 3746
           ,x"8620" -- 3748
           ,x"ed18" -- 374A
           ,x"14f8" -- 374C
           ,x"c818" -- 374E
           ,x"ed18" -- 3750
           ,x"c1e0" -- 3752
           ,x"ed04" -- 3754
           ,x"c078" -- 3756
           ,x"06a0" -- 3758
           ,x"ac2c" -- 375A
           ,x"06a0" -- 375C
           ,x"a37a" -- 375E
           ,x"10eb" -- 3760
           ,x"c2e0" -- 3762
           ,x"ed16" -- 3764
           ,x"045b" -- 3766
           ,x"c032" -- 3768
           ,x"1602" -- 376A
           ,x"c012" -- 376C
           ,x"1306" -- 376E
           ,x"1503" -- 3770
           ,x"0620" -- 3772
           ,x"ef6a" -- 3774
           ,x"1002" -- 3776
           ,x"05a0" -- 3778
           ,x"ef6a" -- 377A
           ,x"0460" -- 377C
           ,x"b6be" -- 377E
           ,x"06a0" -- 3780
           ,x"a226" -- 3782
           ,x"0a0d" -- 3784
           ,x"5052" -- 3786
           ,x"474d" -- 3788
           ,x"c600" -- 378A
           ,x"c060" -- 378C
           ,x"edd8" -- 378E
           ,x"6060" -- 3790
           ,x"edd6" -- 3792
           ,x"a060" -- 3794
           ,x"edd4" -- 3796
           ,x"6060" -- 3798
           ,x"ed0e" -- 379A
           ,x"06a0" -- 379C
           ,x"a1e6" -- 379E
           ,x"06a0" -- 37A0
           ,x"a202" -- 37A2
           ,x"5641" -- 37A4
           ,x"5253" -- 37A6
           ,x"c600" -- 37A8
           ,x"c060" -- 37AA
           ,x"ed04" -- 37AC
           ,x"6060" -- 37AE
           ,x"edda" -- 37B0
           ,x"a060" -- 37B2
           ,x"edd8" -- 37B4
           ,x"6060" -- 37B6
           ,x"edd6" -- 37B8
           ,x"0221" -- 37BA
           ,x"fff8" -- 37BC
           ,x"06a0" -- 37BE
           ,x"a1e6" -- 37C0
           ,x"06a0" -- 37C2
           ,x"a202" -- 37C4
           ,x"4652" -- 37C6
           ,x"4545" -- 37C8
           ,x"c600" -- 37CA
           ,x"c060" -- 37CC
           ,x"edda" -- 37CE
           ,x"6060" -- 37D0
           ,x"edd8" -- 37D2
           ,x"06a0" -- 37D4
           ,x"a1e6" -- 37D6
           ,x"06a0" -- 37D8
           ,x"a202" -- 37DA
           ,x"0000" -- 37DC
           ,x"0420" -- 37DE
           ,x"8190" -- 37E0
           ,x"0460" -- 37E2
           ,x"8124" -- 37E4
           ,x"0200" -- 37E6
           ,x"ef68" -- 37E8
           ,x"cc20" -- 37EA
           ,x"c838" -- 37EC
           ,x"04f0" -- 37EE
           ,x"c401" -- 37F0
           ,x"0420" -- 37F2
           ,x"bd46" -- 37F4
           ,x"c820" -- 37F6
           ,x"8014" -- 37F8
           ,x"ef9e" -- 37FA
           ,x"0420" -- 37FC
           ,x"b05e" -- 37FE
           ,x"045b" -- 3800
           ,x"c04b" -- 3802
           ,x"06a0" -- 3804
           ,x"a22a" -- 3806
           ,x"2042" -- 3808
           ,x"7974" -- 380A
           ,x"6573" -- 380C
           ,x"0df6" -- 380E
           ,x"c2c1" -- 3810
           ,x"100b" -- 3812
           ,x"c1e0" -- 3814
           ,x"ed04" -- 3816
           ,x"ddfb" -- 3818
           ,x"16fe" -- 381A
           ,x"0607" -- 381C
           ,x"058b" -- 381E
           ,x"024b" -- 3820
           ,x"fffe" -- 3822
           ,x"045b" -- 3824
           ,x"c1e0" -- 3826
           ,x"ed04" -- 3828
           ,x"ddfb" -- 382A
           ,x"13f7" -- 382C
           ,x"15fd" -- 382E
           ,x"c80b" -- 3830
           ,x"ed2c" -- 3832
           ,x"04cb" -- 3834
           ,x"d2e7" -- 3836
           ,x"ffff" -- 3838
           ,x"050b" -- 383A
           ,x"d9cb" -- 383C
           ,x"ffff" -- 383E
           ,x"c2e0" -- 3840
           ,x"ed2c" -- 3842
           ,x"10ec" -- 3844
           ,x"0420" -- 3846
           ,x"8d70" -- 3848
           ,x"0032" -- 384A
           ,x"0420" -- 384C
           ,x"8d70" -- 384E
           ,x"0032" -- 3850
           ,x"0720" -- 3852
           ,x"ed30" -- 3854
           ,x"0460" -- 3856
           ,x"aef8" -- 3858
           ,x"04e0" -- 385A
           ,x"ed30" -- 385C
           ,x"10fb" -- 385E
           ,x"c820" -- 3860
           ,x"801a" -- 3862
           ,x"ef9e" -- 3864
           ,x"0420" -- 3866
           ,x"b558" -- 3868
           ,x"0202" -- 386A
           ,x"8044" -- 386C
           ,x"0204" -- 386E
           ,x"e481" -- 3870
           ,x"c001" -- 3872
           ,x"1310" -- 3874
           ,x"0740" -- 3876
           ,x"1502" -- 3878
           ,x"0204" -- 387A
           ,x"4481" -- 387C
           ,x"0201" -- 387E
           ,x"0001" -- 3880
           ,x"0600" -- 3882
           ,x"1304" -- 3884
           ,x"0280" -- 3886
           ,x"0010" -- 3888
           ,x"1407" -- 388A
           ,x"0a01" -- 388C
           ,x"0484" -- 388E
           ,x"0608" -- 3890
           ,x"0460" -- 3892
           ,x"aef8" -- 3894
           ,x"04d2" -- 3896
           ,x"10fb" -- 3898
           ,x"0420" -- 389A
           ,x"8d70" -- 389C
           ,x"002e" -- 389E
           ,x"0420" -- 38A0
           ,x"8d70" -- 38A2
           ,x"0032" -- 38A4
           ,x"c220" -- 38A6
           ,x"edd2" -- 38A8
           ,x"c338" -- 38AA
           ,x"1305" -- 38AC
           ,x"804c" -- 38AE
           ,x"1302" -- 38B0
           ,x"05c8" -- 38B2
           ,x"10fa" -- 38B4
           ,x"045b" -- 38B6
           ,x"0420" -- 38B8
           ,x"8d70" -- 38BA
           ,x"000d" -- 38BC
           ,x"c020" -- 38BE
           ,x"804c" -- 38C0
           ,x"1602" -- 38C2
           ,x"0460" -- 38C4
           ,x"a36e" -- 38C6
           ,x"c048" -- 38C8
           ,x"0208" -- 38CA
           ,x"2000" -- 38CC
           ,x"0202" -- 38CE
           ,x"1800" -- 38D0
           ,x"06a0" -- 38D2
           ,x"8444" -- 38D4
           ,x"0588" -- 38D6
           ,x"d0e0" -- 38D8
           ,x"0000" -- 38DA
           ,x"c143" -- 38DC
           ,x"0983" -- 38DE
           ,x"c103" -- 38E0
           ,x"0243" -- 38E2
           ,x"000f" -- 38E4
           ,x"d023" -- 38E6
           ,x"8084" -- 38E8
           ,x"0940" -- 38EA
           ,x"0944" -- 38EC
           ,x"d024" -- 38EE
           ,x"8084" -- 38F0
           ,x"0a40" -- 38F2
           ,x"9140" -- 38F4
           ,x"1308" -- 38F6
           ,x"0228" -- 38F8
           ,x"3fff" -- 38FA
           ,x"06a0" -- 38FC
           ,x"8444" -- 38FE
           ,x"0228" -- 3900
           ,x"c001" -- 3902
           ,x"d800" -- 3904
           ,x"0000" -- 3906
           ,x"0602" -- 3908
           ,x"16e3" -- 390A
           ,x"c201" -- 390C
           ,x"0460" -- 390E
           ,x"aef8" -- 3910
           ,x"0420" -- 3912
           ,x"be74" -- 3914
           ,x"c0f1" -- 3916
           ,x"1602" -- 3918
           ,x"c0d1" -- 391A
           ,x"1306" -- 391C
           ,x"c0f2" -- 391E
           ,x"1602" -- 3920
           ,x"c0d2" -- 3922
           ,x"1302" -- 3924
           ,x"05a0" -- 3926
           ,x"ef6a" -- 3928
           ,x"0202" -- 392A
           ,x"ef68" -- 392C
           ,x"045b" -- 392E
           ,x"0420" -- 3930
           ,x"be74" -- 3932
           ,x"c0f1" -- 3934
           ,x"16f7" -- 3936
           ,x"c0d1" -- 3938
           ,x"16f5" -- 393A
           ,x"c0f2" -- 393C
           ,x"16f3" -- 393E
           ,x"c0d2" -- 3940
           ,x"16f1" -- 3942
           ,x"10f2" -- 3944
           ,x"0420" -- 3946
           ,x"be74" -- 3948
           ,x"c0f1" -- 394A
           ,x"16ee" -- 394C
           ,x"c0d1" -- 394E
           ,x"13ea" -- 3950
           ,x"10eb" -- 3952
           ,x"0720" -- 3954
           ,x"ede4" -- 3956
           ,x"0420" -- 3958
           ,x"8170" -- 395A
           ,x"c060" -- 395C
           ,x"ed32" -- 395E
           ,x"0460" -- 3960
           ,x"9502" -- 3962
           ,x"c820" -- 3964
           ,x"ede4" -- 3966
           ,x"ede4" -- 3968
           ,x"1601" -- 396A
           ,x"045b" -- 396C
           ,x"0420" -- 396E
           ,x"8d70" -- 3970
           ,x"0030" -- 3972
           ,x"c820" -- 3974
           ,x"9f86" -- 3976
           ,x"ed14" -- 3978
           ,x"c28b" -- 397A
           ,x"c806" -- 397C
           ,x"ed02" -- 397E
           ,x"04e0" -- 3980
           ,x"8042" -- 3982
           ,x"c1e0" -- 3984
           ,x"ed04" -- 3986
           ,x"0206" -- 3988
           ,x"ee82" -- 398A
           ,x"0716" -- 398C
           ,x"0208" -- 398E
           ,x"edfe" -- 3990
           ,x"c160" -- 3992
           ,x"edd4" -- 3994
           ,x"04f5" -- 3996
           ,x"04f5" -- 3998
           ,x"04f5" -- 399A
           ,x"0200" -- 399C
           ,x"11d2" -- 399E
           ,x"c540" -- 39A0
           ,x"0420" -- 39A2
           ,x"b284" -- 39A4
           ,x"1042" -- 39A6
           ,x"04c1" -- 39A8
           ,x"c801" -- 39AA
           ,x"edee" -- 39AC
           ,x"113e" -- 39AE
           ,x"1301" -- 39B0
           ,x"0607" -- 39B2
           ,x"c000" -- 39B4
           ,x"1608" -- 39B6
           ,x"c2e0" -- 39B8
           ,x"ede0" -- 39BA
           ,x"1602" -- 39BC
           ,x"0460" -- 39BE
           ,x"a77e" -- 39C0
           ,x"04e0" -- 39C2
           ,x"ede0" -- 39C4
           ,x"045a" -- 39C6
           ,x"06a0" -- 39C8
           ,x"a92c" -- 39CA
           ,x"1038" -- 39CC
           ,x"c0c7" -- 39CE
           ,x"c001" -- 39D0
           ,x"06a0" -- 39D2
           ,x"a934" -- 39D4
           ,x"1014" -- 39D6
           ,x"a001" -- 39D8
           ,x"0280" -- 39DA
           ,x"1920" -- 39DC
           ,x"1329" -- 39DE
           ,x"0280" -- 39E0
           ,x"39e0" -- 39E2
           ,x"1329" -- 39E4
           ,x"06a0" -- 39E6
           ,x"a934" -- 39E8
           ,x"100a" -- 39EA
           ,x"a001" -- 39EC
           ,x"0204" -- 39EE
           ,x"a99c" -- 39F0
           ,x"c074" -- 39F2
           ,x"0911" -- 39F4
           ,x"8040" -- 39F6
           ,x"1307" -- 39F8
           ,x"0284" -- 39FA
           ,x"aa48" -- 39FC
           ,x"1af9" -- 39FE
           ,x"c1c3" -- 3A00
           ,x"de20" -- 3A02
           ,x"ac6e" -- 3A04
           ,x"105c" -- 3A06
           ,x"c080" -- 3A08
           ,x"c3c7" -- 3A0A
           ,x"c024" -- 3A0C
           ,x"00aa" -- 3A0E
           ,x"1733" -- 3A10
           ,x"c140" -- 3A12
           ,x"0245" -- 3A14
           ,x"003e" -- 3A16
           ,x"132f" -- 3A18
           ,x"06a0" -- 3A1A
           ,x"a934" -- 3A1C
           ,x"1003" -- 3A1E
           ,x"0991" -- 3A20
           ,x"8045" -- 3A22
           ,x"13f6" -- 3A24
           ,x"c002" -- 3A26
           ,x"c1cf" -- 3A28
           ,x"10e3" -- 3A2A
           ,x"06a0" -- 3A2C
           ,x"c0f6" -- 3A2E
           ,x"3033" -- 3A30
           ,x"0204" -- 3A32
           ,x"0082" -- 3A34
           ,x"102a" -- 3A36
           ,x"0204" -- 3A38
           ,x"0080" -- 3A3A
           ,x"1027" -- 3A3C
           ,x"9817" -- 3A3E
           ,x"c8d6" -- 3A40
           ,x"160d" -- 3A42
           ,x"0587" -- 3A44
           ,x"0204" -- 3A46
           ,x"4600" -- 3A48
           ,x"de04" -- 3A4A
           ,x"d037" -- 3A4C
           ,x"1305" -- 3A4E
           ,x"9800" -- 3A50
           ,x"c0e4" -- 3A52
           ,x"1302" -- 3A54
           ,x"de00" -- 3A56
           ,x"10f9" -- 3A58
           ,x"7e18" -- 3A5A
           ,x"1032" -- 3A5C
           ,x"9837" -- 3A5E
           ,x"c8c0" -- 3A60
           ,x"1603" -- 3A62
           ,x"0204" -- 3A64
           ,x"008a" -- 3A66
           ,x"1011" -- 3A68
           ,x"0607" -- 3A6A
           ,x"9837" -- 3A6C
           ,x"ab6d" -- 3A6E
           ,x"16c8" -- 3A70
           ,x"0204" -- 3A72
           ,x"007e" -- 3A74
           ,x"100a" -- 3A76
           ,x"0201" -- 3A78
           ,x"a9b2" -- 3A7A
           ,x"6101" -- 3A7C
           ,x"1506" -- 3A7E
           ,x"c000" -- 3A80
           ,x"1301" -- 3A82
           ,x"0450" -- 3A84
           ,x"0420" -- 3A86
           ,x"8d70" -- 3A88
           ,x"ffff" -- 3A8A
           ,x"e820" -- 3A8C
           ,x"b920" -- 3A8E
           ,x"8046" -- 3A90
           ,x"0a74" -- 3A92
           ,x"de04" -- 3A94
           ,x"0284" -- 3A96
           ,x"0300" -- 3A98
           ,x"1108" -- 3A9A
           ,x"1395" -- 3A9C
           ,x"0284" -- 3A9E
           ,x"0400" -- 3AA0
           ,x"160f" -- 3AA2
           ,x"0460" -- 3AA4
           ,x"a6c0" -- 3AA6
           ,x"de20" -- 3AA8
           ,x"c8c0" -- 3AAA
           ,x"0420" -- 3AAC
           ,x"b284" -- 3AAE
           ,x"1000" -- 3AB0
           ,x"10bc" -- 3AB2
           ,x"de01" -- 3AB4
           ,x"06c1" -- 3AB6
           ,x"de01" -- 3AB8
           ,x"0280" -- 3ABA
           ,x"2c00" -- 3ABC
           ,x"13f4" -- 3ABE
           ,x"0607" -- 3AC0
           ,x"c308" -- 3AC2
           ,x"0420" -- 3AC4
           ,x"b288" -- 3AC6
           ,x"1014" -- 3AC8
           ,x"101d" -- 3ACA
           ,x"1009" -- 3ACC
           ,x"0281" -- 3ACE
           ,x"ffff" -- 3AD0
           ,x"1109" -- 3AD2
           ,x"8801" -- 3AD4
           ,x"ed14" -- 3AD6
           ,x"1506" -- 3AD8
           ,x"0221" -- 3ADA
           ,x"0063" -- 3ADC
           ,x"1006" -- 3ADE
           ,x"de20" -- 3AE0
           ,x"adeb" -- 3AE2
           ,x"1002" -- 3AE4
           ,x"de20" -- 3AE6
           ,x"ab7c" -- 3AE8
           ,x"de01" -- 3AEA
           ,x"06c1" -- 3AEC
           ,x"de01" -- 3AEE
           ,x"1009" -- 3AF0
           ,x"de20" -- 3AF2
           ,x"ab7e" -- 3AF4
           ,x"0203" -- 3AF6
           ,x"0006" -- 3AF8
           ,x"0204" -- 3AFA
           ,x"ef68" -- 3AFC
           ,x"de34" -- 3AFE
           ,x"0603" -- 3B00
           ,x"16fd" -- 3B02
           ,x"0607" -- 3B04
           ,x"06a0" -- 3B06
           ,x"a94c" -- 3B08
           ,x"06a0" -- 3B0A
           ,x"a92c" -- 3B0C
           ,x"1062" -- 3B0E
           ,x"c001" -- 3B10
           ,x"06a0" -- 3B12
           ,x"a934" -- 3B14
           ,x"101d" -- 3B16
           ,x"a001" -- 3B18
           ,x"0280" -- 3B1A
           ,x"38c0" -- 3B1C
           ,x"1602" -- 3B1E
           ,x"0460" -- 3B20
           ,x"a70c" -- 3B22
           ,x"06a0" -- 3B24
           ,x"a934" -- 3B26
           ,x"1025" -- 3B28
           ,x"a001" -- 3B2A
           ,x"0204" -- 3B2C
           ,x"aace" -- 3B2E
           ,x"c074" -- 3B30
           ,x"0911" -- 3B32
           ,x"8040" -- 3B34
           ,x"1609" -- 3B36
           ,x"020b" -- 3B38
           ,x"aace" -- 3B3A
           ,x"0224" -- 3B3C
           ,x"0034" -- 3B3E
           ,x"610b" -- 3B40
           ,x"0914" -- 3B42
           ,x"06c4" -- 3B44
           ,x"de04" -- 3B46
           ,x"10bd" -- 3B48
           ,x"0284" -- 3B4A
           ,x"ab08" -- 3B4C
           ,x"1af0" -- 3B4E
           ,x"1011" -- 3B50
           ,x"c0c0" -- 3B52
           ,x"06a0" -- 3B54
           ,x"b416" -- 3B56
           ,x"100b" -- 3B58
           ,x"0607" -- 3B5A
           ,x"0420" -- 3B5C
           ,x"b284" -- 3B5E
           ,x"101f" -- 3B60
           ,x"1007" -- 3B62
           ,x"2460" -- 3B64
           ,x"aa66" -- 3B66
           ,x"161b" -- 3B68
           ,x"a0c1" -- 3B6A
           ,x"0263" -- 3B6C
           ,x"0380" -- 3B6E
           ,x"0607" -- 3B70
           ,x"c003" -- 3B72
           ,x"06a0" -- 3B74
           ,x"a982" -- 3B76
           ,x"1002" -- 3B78
           ,x"0607" -- 3B7A
           ,x"1003" -- 3B7C
           ,x"0500" -- 3B7E
           ,x"05c6" -- 3B80
           ,x"0716" -- 3B82
           ,x"0204" -- 3B84
           ,x"ff70" -- 3B86
           ,x"c160" -- 3B88
           ,x"edd4" -- 3B8A
           ,x"8805" -- 3B8C
           ,x"edd6" -- 3B8E
           ,x"140d" -- 3B90
           ,x"8d40" -- 3B92
           ,x"131b" -- 3B94
           ,x"0584" -- 3B96
           ,x"16f9" -- 3B98
           ,x"0420" -- 3B9A
           ,x"8d70" -- 3B9C
           ,x"0005" -- 3B9E
           ,x"06a0" -- 3BA0
           ,x"c0f6" -- 3BA2
           ,x"3034" -- 3BA4
           ,x"0420" -- 3BA6
           ,x"8d70" -- 3BA8
           ,x"000a" -- 3BAA
           ,x"c0a0" -- 3BAC
           ,x"edd8" -- 3BAE
           ,x"8cb2" -- 3BB0
           ,x"8802" -- 3BB2
           ,x"edda" -- 3BB4
           ,x"14f7" -- 3BB6
           ,x"c802" -- 3BB8
           ,x"edd8" -- 3BBA
           ,x"0222" -- 3BBC
           ,x"fffc" -- 3BBE
           ,x"c4b2" -- 3BC0
           ,x"8142" -- 3BC2
           ,x"1bfb" -- 3BC4
           ,x"c540" -- 3BC6
           ,x"05e0" -- 3BC8
           ,x"edd6" -- 3BCA
           ,x"c000" -- 3BCC
           ,x"11ba" -- 3BCE
           ,x"06c4" -- 3BD0
           ,x"de04" -- 3BD2
           ,x"04c0" -- 3BD4
           ,x"d037" -- 3BD6
           ,x"1375" -- 3BD8
           ,x"c040" -- 3BDA
           ,x"06c1" -- 3BDC
           ,x"0280" -- 3BDE
           ,x"4100" -- 3BE0
           ,x"1a08" -- 3BE2
           ,x"0280" -- 3BE4
           ,x"5b00" -- 3BE6
           ,x"1a47" -- 3BE8
           ,x"0221" -- 3BEA
           ,x"ffe6" -- 3BEC
           ,x"0280" -- 3BEE
           ,x"5e00" -- 3BF0
           ,x"1b3f" -- 3BF2
           ,x"d061" -- 3BF4
           ,x"aae9" -- 3BF6
           ,x"133c" -- 3BF8
           ,x"d601" -- 3BFA
           ,x"06a0" -- 3BFC
           ,x"872c" -- 3BFE
           ,x"ea20" -- 3C00
           ,x"4228" -- 3C02
           ,x"425b" -- 3C04
           ,x"5529" -- 3C06
           ,x"555d" -- 3C08
           ,x"0f22" -- 3C0A
           ,x"0f27" -- 3C0C
           ,x"303a" -- 3C0E
           ,x"5f21" -- 3C10
           ,x"163d" -- 3C12
           ,x"273e" -- 3C14
           ,x"0000" -- 3C16
           ,x"0588" -- 3C18
           ,x"0460" -- 3C1A
           ,x"a4c4" -- 3C1C
           ,x"0588" -- 3C1E
           ,x"d637" -- 3C20
           ,x"1371" -- 3C22
           ,x"9600" -- 3C24
           ,x"16fb" -- 3C26
           ,x"7e18" -- 3C28
           ,x"10f7" -- 3C2A
           ,x"0608" -- 3C2C
           ,x"9818" -- 3C2E
           ,x"ab27" -- 3C30
           ,x"130a" -- 3C32
           ,x"9818" -- 3C34
           ,x"ab25" -- 3C36
           ,x"1307" -- 3C38
           ,x"9838" -- 3C3A
           ,x"ab26" -- 3C3C
           ,x"16ec" -- 3C3E
           ,x"7a20" -- 3C40
           ,x"b921" -- 3C42
           ,x"ffff" -- 3C44
           ,x"10e9" -- 3C46
           ,x"be20" -- 3C48
           ,x"b921" -- 3C4A
           ,x"10e6" -- 3C4C
           ,x"9828" -- 3C4E
           ,x"ffff" -- 3C50
           ,x"ab25" -- 3C52
           ,x"16e1" -- 3C54
           ,x"ba20" -- 3C56
           ,x"aa6b" -- 3C58
           ,x"ffff" -- 3C5A
           ,x"10de" -- 3C5C
           ,x"0587" -- 3C5E
           ,x"9817" -- 3C60
           ,x"c0e4" -- 3C62
           ,x"13fc" -- 3C64
           ,x"9817" -- 3C66
           ,x"c8dd" -- 3C68
           ,x"13f9" -- 3C6A
           ,x"0588" -- 3C6C
           ,x"0460" -- 3C6E
           ,x"a3c8" -- 3C70
           ,x"06a0" -- 3C72
           ,x"c0f6" -- 3C74
           ,x"3036" -- 3C76
           ,x"0607" -- 3C78
           ,x"06a0" -- 3C7A
           ,x"a94c" -- 3C7C
           ,x"06a0" -- 3C7E
           ,x"c0f6" -- 3C80
           ,x"3037" -- 3C82
           ,x"8308" -- 3C84
           ,x"1b05" -- 3C86
           ,x"9828" -- 3C88
           ,x"ffff" -- 3C8A
           ,x"aa64" -- 3C8C
           ,x"1a0b" -- 3C8E
           ,x"1006" -- 3C90
           ,x"d068" -- 3C92
           ,x"ffff" -- 3C94
           ,x"1307" -- 3C96
           ,x"9801" -- 3C98
           ,x"ab7f" -- 3C9A
           ,x"1404" -- 3C9C
           ,x"05c6" -- 3C9E
           ,x"04d6" -- 3CA0
           ,x"7620" -- 3CA2
           ,x"aa6b" -- 3CA4
           ,x"0616" -- 3CA6
           ,x"10b7" -- 3CA8
           ,x"0596" -- 3CAA
           ,x"1106" -- 3CAC
           ,x"0646" -- 3CAE
           ,x"0286" -- 3CB0
           ,x"ee82" -- 3CB2
           ,x"1a28" -- 3CB4
           ,x"7620" -- 3CB6
           ,x"aa6b" -- 3CB8
           ,x"0588" -- 3CBA
           ,x"108b" -- 3CBC
           ,x"0588" -- 3CBE
           ,x"de37" -- 3CC0
           ,x"16fe" -- 3CC2
           ,x"0286" -- 3CC4
           ,x"ee82" -- 3CC6
           ,x"161e" -- 3CC8
           ,x"0596" -- 3CCA
           ,x"161c" -- 3CCC
           ,x"7e18" -- 3CCE
           ,x"7618" -- 3CD0
           ,x"0700" -- 3CD2
           ,x"c060" -- 3CD4
           ,x"edee" -- 3CD6
           ,x"1652" -- 3CD8
           ,x"c1e0" -- 3CDA
           ,x"ed04" -- 3CDC
           ,x"0227" -- 3CDE
           ,x"001e" -- 3CE0
           ,x"c007" -- 3CE2
           ,x"0203" -- 3CE4
           ,x"edfe" -- 3CE6
           ,x"cdf3" -- 3CE8
           ,x"8203" -- 3CEA
           ,x"1afd" -- 3CEC
           ,x"04e0" -- 3CEE
           ,x"8046" -- 3CF0
           ,x"c200" -- 3CF2
           ,x"9818" -- 3CF4
           ,x"b921" -- 3CF6
           ,x"1b04" -- 3CF8
           ,x"0720" -- 3CFA
           ,x"ede4" -- 3CFC
           ,x"0420" -- 3CFE
           ,x"8170" -- 3D00
           ,x"0460" -- 3D02
           ,x"af38" -- 3D04
           ,x"06a0" -- 3D06
           ,x"c0f6" -- 3D08
           ,x"3032" -- 3D0A
           ,x"06a0" -- 3D0C
           ,x"a92c" -- 3D0E
           ,x"102f" -- 3D10
           ,x"0921" -- 3D12
           ,x"de01" -- 3D14
           ,x"c0c8" -- 3D16
           ,x"0643" -- 3D18
           ,x"0283" -- 3D1A
           ,x"edfe" -- 3D1C
           ,x"16ce" -- 3D1E
           ,x"9813" -- 3D20
           ,x"ab80" -- 3D22
           ,x"16cb" -- 3D24
           ,x"06a0" -- 3D26
           ,x"a982" -- 3D28
           ,x"1002" -- 3D2A
           ,x"0607" -- 3D2C
           ,x"1017" -- 3D2E
           ,x"0203" -- 3D30
           ,x"0003" -- 3D32
           ,x"c120" -- 3D34
           ,x"edd4" -- 3D36
           ,x"06a0" -- 3D38
           ,x"a92c" -- 3D3A
           ,x"101c" -- 3D3C
           ,x"de01" -- 3D3E
           ,x"cd01" -- 3D40
           ,x"06a0" -- 3D42
           ,x"a982" -- 3D44
           ,x"1017" -- 3D46
           ,x"0603" -- 3D48
           ,x"1303" -- 3D4A
           ,x"0281" -- 3D4C
           ,x"2c00" -- 3D4E
           ,x"13f3" -- 3D50
           ,x"0281" -- 3D52
           ,x"2900" -- 3D54
           ,x"1303" -- 3D56
           ,x"0281" -- 3D58
           ,x"5d00" -- 3D5A
           ,x"16d4" -- 3D5C
           ,x"95e0" -- 3D5E
           ,x"ab83" -- 3D60
           ,x"13ac" -- 3D62
           ,x"9de0" -- 3D64
           ,x"c0e4" -- 3D66
           ,x"13fa" -- 3D68
           ,x"06a0" -- 3D6A
           ,x"c0f6" -- 3D6C
           ,x"3336" -- 3D6E
           ,x"06a0" -- 3D70
           ,x"c0f6" -- 3D72
           ,x"3038" -- 3D74
           ,x"06a0" -- 3D76
           ,x"c0f6" -- 3D78
           ,x"3039" -- 3D7A
           ,x"c28b" -- 3D7C
           ,x"c041" -- 3D7E
           ,x"1377" -- 3D80
           ,x"0202" -- 3D82
           ,x"edfe" -- 3D84
           ,x"6202" -- 3D86
           ,x"0588" -- 3D88
           ,x"0818" -- 3D8A
           ,x"c088" -- 3D8C
           ,x"a082" -- 3D8E
           ,x"c1a0" -- 3D90
           ,x"edd2" -- 3D92
           ,x"c1c6" -- 3D94
           ,x"61e0" -- 3D96
           ,x"ed0e" -- 3D98
           ,x"c116" -- 3D9A
           ,x"1309" -- 3D9C
           ,x"8581" -- 3D9E
           ,x"1368" -- 3DA0
           ,x"1506" -- 3DA2
           ,x"05c6" -- 3DA4
           ,x"c1f6" -- 3DA6
           ,x"10f8" -- 3DA8
           ,x"0420" -- 3DAA
           ,x"8d70" -- 3DAC
           ,x"000d" -- 3DAE
           ,x"c000" -- 3DB0
           ,x"13fb" -- 3DB2
           ,x"c0c6" -- 3DB4
           ,x"06a0" -- 3DB6
           ,x"a8aa" -- 3DB8
           ,x"0004" -- 3DBA
           ,x"cd81" -- 3DBC
           ,x"c587" -- 3DBE
           ,x"0204" -- 3DC0
           ,x"edfe" -- 3DC2
           ,x"c196" -- 3DC4
           ,x"a1a0" -- 3DC6
           ,x"ed0e" -- 3DC8
           ,x"c1c6" -- 3DCA
           ,x"cdf4" -- 3DCC
           ,x"0608" -- 3DCE
           ,x"16fd" -- 3DD0
           ,x"c120" -- 3DD2
           ,x"eddc" -- 3DD4
           ,x"8804" -- 3DD6
           ,x"ed0a" -- 3DD8
           ,x"1217" -- 3DDA
           ,x"0224" -- 3DDC
           ,x"fffc" -- 3DDE
           ,x"8506" -- 3DE0
           ,x"1b0e" -- 3DE2
           ,x"8507" -- 3DE4
           ,x"120a" -- 3DE6
           ,x"c144" -- 3DE8
           ,x"cd65" -- 3DEA
           ,x"0004" -- 3DEC
           ,x"8805" -- 3DEE
           ,x"eddc" -- 3DF0
           ,x"1afb" -- 3DF2
           ,x"a820" -- 3DF4
           ,x"a886" -- 3DF6
           ,x"eddc" -- 3DF8
           ,x"10ed" -- 3DFA
           ,x"a502" -- 3DFC
           ,x"1002" -- 3DFE
           ,x"a903" -- 3E00
           ,x"0002" -- 3E02
           ,x"a902" -- 3E04
           ,x"0002" -- 3E06
           ,x"10e6" -- 3E08
           ,x"c120" -- 3E0A
           ,x"ed08" -- 3E0C
           ,x"c014" -- 3E0E
           ,x"1313" -- 3E10
           ,x"c144" -- 3E12
           ,x"0225" -- 3E14
           ,x"000e" -- 3E16
           ,x"8546" -- 3E18
           ,x"1b07" -- 3E1A
           ,x"8547" -- 3E1C
           ,x"1203" -- 3E1E
           ,x"06a0" -- 3E20
           ,x"9142" -- 3E22
           ,x"10f4" -- 3E24
           ,x"a542" -- 3E26
           ,x"1002" -- 3E28
           ,x"a943" -- 3E2A
           ,x"0002" -- 3E2C
           ,x"a942" -- 3E2E
           ,x"0002" -- 3E30
           ,x"0224" -- 3E32
           ,x"0012" -- 3E34
           ,x"10eb" -- 3E36
           ,x"0204" -- 3E38
           ,x"edec" -- 3E3A
           ,x"8506" -- 3E3C
           ,x"1b09" -- 3E3E
           ,x"8507" -- 3E40
           ,x"1202" -- 3E42
           ,x"04d4" -- 3E44
           ,x"1003" -- 3E46
           ,x"c014" -- 3E48
           ,x"1303" -- 3E4A
           ,x"a502" -- 3E4C
           ,x"a803" -- 3E4E
           ,x"edea" -- 3E50
           ,x"c120" -- 3E52
           ,x"ed0c" -- 3E54
           ,x"c014" -- 3E56
           ,x"1307" -- 3E58
           ,x"8506" -- 3E5A
           ,x"1b05" -- 3E5C
           ,x"8507" -- 3E5E
           ,x"1202" -- 3E60
           ,x"04d4" -- 3E62
           ,x"1001" -- 3E64
           ,x"a502" -- 3E66
           ,x"8d34" -- 3E68
           ,x"8804" -- 3E6A
           ,x"ed0a" -- 3E6C
           ,x"1af3" -- 3E6E
           ,x"045a" -- 3E70
           ,x"c2e6" -- 3E72
           ,x"0002" -- 3E74
           ,x"62c7" -- 3E76
           ,x"c000" -- 3E78
           ,x"1607" -- 3E7A
           ,x"c08b" -- 3E7C
           ,x"c0c6" -- 3E7E
           ,x"8cf3" -- 3E80
           ,x"06a0" -- 3E82
           ,x"a8aa" -- 3E84
           ,x"fffc" -- 3E86
           ,x"10a4" -- 3E88
           ,x"a08b" -- 3E8A
           ,x"c020" -- 3E8C
           ,x"edd8" -- 3E8E
           ,x"a002" -- 3E90
           ,x"8800" -- 3E92
           ,x"edda" -- 3E94
           ,x"1406" -- 3E96
           ,x"020d" -- 3E98
           ,x"a89e" -- 3E9A
           ,x"1019" -- 3E9C
           ,x"0000" -- 3E9E
           ,x"05c6" -- 3EA0
           ,x"108e" -- 3EA2
           ,x"0420" -- 3EA4
           ,x"8d70" -- 3EA6
           ,x"000a" -- 3EA8
           ,x"c34b" -- 3EAA
           ,x"c120" -- 3EAC
           ,x"edd8" -- 3EAE
           ,x"c143" -- 3EB0
           ,x"a15d" -- 3EB2
           ,x"c004" -- 3EB4
           ,x"a01d" -- 3EB6
           ,x"a002" -- 3EB8
           ,x"8800" -- 3EBA
           ,x"edda" -- 3EBC
           ,x"14f2" -- 3EBE
           ,x"a81d" -- 3EC0
           ,x"edd4" -- 3EC2
           ,x"a81d" -- 3EC4
           ,x"edd6" -- 3EC6
           ,x"a81d" -- 3EC8
           ,x"edd8" -- 3ECA
           ,x"06a0" -- 3ECC
           ,x"a90c" -- 3ECE
           ,x"c0c7" -- 3ED0
           ,x"a0e0" -- 3ED2
           ,x"ed0e" -- 3ED4
           ,x"c120" -- 3ED6
           ,x"edd8" -- 3ED8
           ,x"c143" -- 3EDA
           ,x"a142" -- 3EDC
           ,x"a182" -- 3EDE
           ,x"a802" -- 3EE0
           ,x"edd2" -- 3EE2
           ,x"a802" -- 3EE4
           ,x"edd4" -- 3EE6
           ,x"a802" -- 3EE8
           ,x"edd6" -- 3EEA
           ,x"a802" -- 3EEC
           ,x"edd8" -- 3EEE
           ,x"a802" -- 3EF0
           ,x"ed2a" -- 3EF2
           ,x"06a0" -- 3EF4
           ,x"a90c" -- 3EF6
           ,x"c0c6" -- 3EF8
           ,x"8803" -- 3EFA
           ,x"edd2" -- 3EFC
           ,x"1204" -- 3EFE
           ,x"0643" -- 3F00
           ,x"a4c2" -- 3F02
           ,x"0643" -- 3F04
           ,x"10f9" -- 3F06
           ,x"c0fd" -- 3F08
           ,x"045d" -- 3F0A
           ,x"8143" -- 3F0C
           ,x"131d" -- 3F0E
           ,x"1a04" -- 3F10
           ,x"8103" -- 3F12
           ,x"1b1a" -- 3F14
           ,x"cd73" -- 3F16
           ,x"10fc" -- 3F18
           ,x"c004" -- 3F1A
           ,x"6003" -- 3F1C
           ,x"a140" -- 3F1E
           ,x"c554" -- 3F20
           ,x"8103" -- 3F22
           ,x"1312" -- 3F24
           ,x"0644" -- 3F26
           ,x"0645" -- 3F28
           ,x"10fa" -- 3F2A
           ,x"9de0" -- 3F2C
           ,x"c0e4" -- 3F2E
           ,x"13fd" -- 3F30
           ,x"0607" -- 3F32
           ,x"9817" -- 3F34
           ,x"c8e0" -- 3F36
           ,x"1208" -- 3F38
           ,x"9817" -- 3F3A
           ,x"ab77" -- 3F3C
           ,x"1405" -- 3F3E
           ,x"04c1" -- 3F40
           ,x"d077" -- 3F42
           ,x"0a21" -- 3F44
           ,x"0950" -- 3F46
           ,x"05cb" -- 3F48
           ,x"045b" -- 3F4A
           ,x"c14b" -- 3F4C
           ,x"06a0" -- 3F4E
           ,x"a92c" -- 3F50
           ,x"0455" -- 3F52
           ,x"0607" -- 3F54
           ,x"0204" -- 3F56
           ,x"ab2e" -- 3F58
           ,x"c0c7" -- 3F5A
           ,x"d074" -- 3F5C
           ,x"1308" -- 3F5E
           ,x"9073" -- 3F60
           ,x"13fc" -- 3F62
           ,x"d074" -- 3F64
           ,x"16fe" -- 3F66
           ,x"0584" -- 3F68
           ,x"d054" -- 3F6A
           ,x"16f6" -- 3F6C
           ,x"0455" -- 3F6E
           ,x"d614" -- 3F70
           ,x"c1c3" -- 3F72
           ,x"9818" -- 3F74
           ,x"ab6d" -- 3F76
           ,x"1302" -- 3F78
           ,x"0460" -- 3F7A
           ,x"a618" -- 3F7C
           ,x"0460" -- 3F7E
           ,x"a660" -- 3F80
           ,x"04c1" -- 3F82
           ,x"d077" -- 3F84
           ,x"0281" -- 3F86
           ,x"2000" -- 3F88
           ,x"13fb" -- 3F8A
           ,x"0281" -- 3F8C
           ,x"2800" -- 3F8E
           ,x"1304" -- 3F90
           ,x"0281" -- 3F92
           ,x"5b00" -- 3F94
           ,x"1301" -- 3F96
           ,x"05cb" -- 3F98
           ,x"045b" -- 3F9A
           ,x"7564" -- 3F9C
           ,x"d266" -- 3F9E
           ,x"73c6" -- 3FA0
           ,x"73da" -- 3FA2
           ,x"0000" -- 3FA4
           ,x"0000" -- 3FA6
           ,x"0000" -- 3FA8
           ,x"0000" -- 3FAA
           ,x"0000" -- 3FAC
           ,x"0000" -- 3FAE
           ,x"0000" -- 3FB0
           ,x"a3cf" -- 3FB2
           ,x"9bcf" -- 3FB4
           ,x"9b0b" -- 3FB6
           ,x"6964" -- 3FB8
           ,x"93cc" -- 3FBA
           ,x"0000" -- 3FBC
           ,x"a049" -- 3FBE
           ,x"c15d" -- 3FC0
           ,x"948b" -- 3FC2
           ,x"4ca1" -- 3FC4
           ,x"6047" -- 3FC6
           ,x"0bd9" -- 3FC8
           ,x"8393" -- 3FCA
           ,x"0965" -- 3FCC
           ,x"9965" -- 3FCE
           ,x"a165" -- 3FD0
           ,x"7d27" -- 3FD2
           ,x"4bab" -- 3FD4
           ,x"6a69" -- 3FD6
           ,x"b067" -- 3FD8
           ,x"9845" -- 3FDA
           ,x"1ccb" -- 3FDC
           ,x"2bdd" -- 3FDE
           ,x"7065" -- 3FE0
           ,x"a845" -- 3FE2
           ,x"a38b" -- 3FE4
           ,x"7b21" -- 3FE6
           ,x"83ab" -- 3FE8
           ,x"63c7" -- 3FEA
           ,x"9561" -- 3FEC
           ,x"0c8f" -- 3FEE
           ,x"c169" -- 3FF0
           ,x"486f" -- 3FF2
           ,x"0a07" -- 3FF4
           ,x"6d5d" -- 3FF6
           ,x"9a59" -- 3FF8
           ,x"7165" -- 3FFA
           ,x"9427" -- 3FFC
           ,x"0a27" -- 3FFE
           ,x"ac27" -- 4000
           ,x"29e7" -- 4002
           ,x"7bc5" -- 4004
           ,x"0de7" -- 4006
           ,x"0000" -- 4008
           ,x"a3db" -- 400A
           ,x"0000" -- 400C
           ,x"0000" -- 400E
           ,x"0000" -- 4010
           ,x"0000" -- 4012
           ,x"0000" -- 4014
           ,x"0000" -- 4016
           ,x"0000" -- 4018
           ,x"0000" -- 401A
           ,x"0000" -- 401C
           ,x"0000" -- 401E
           ,x"0000" -- 4020
           ,x"385a" -- 4022
           ,x"33e8" -- 4024
           ,x"73e8" -- 4026
           ,x"83e0" -- 4028
           ,x"6a48" -- 402A
           ,x"a158" -- 402C
           ,x"0000" -- 402E
           ,x"73c0" -- 4030
           ,x"3240" -- 4032
           ,x"3148" -- 4034
           ,x"b95c" -- 4036
           ,x"238a" -- 4038
           ,x"0000" -- 403A
           ,x"0000" -- 403C
           ,x"a244" -- 403E
           ,x"1486" -- 4040
           ,x"3486" -- 4042
           ,x"695a" -- 4044
           ,x"25da" -- 4046
           ,x"aebe" -- 4048
           ,x"a180" -- 404A
           ,x"a354" -- 404C
           ,x"871e" -- 404E
           ,x"0000" -- 4050
           ,x"0000" -- 4052
           ,x"0000" -- 4054
           ,x"0000" -- 4056
           ,x"0000" -- 4058
           ,x"0000" -- 405A
           ,x"0000" -- 405C
           ,x"001e" -- 405E
           ,x"00aa" -- 4060
           ,x"000a" -- 4062
           ,x"4700" -- 4064
           ,x"ff80" -- 4066
           ,x"0000" -- 4068
           ,x"0002" -- 406A
           ,x"0028" -- 406C
           ,x"049e" -- 406E
           ,x"051c" -- 4070
           ,x"0018" -- 4072
           ,x"0008" -- 4074
           ,x"052a" -- 4076
           ,x"0008" -- 4078
           ,x"93e8" -- 407A
           ,x"74aa" -- 407C
           ,x"0020" -- 407E
           ,x"0028" -- 4080
           ,x"000a" -- 4082
           ,x"000a" -- 4084
           ,x"000a" -- 4086
           ,x"2c02" -- 4088
           ,x"00e6" -- 408A
           ,x"6bc8" -- 408C
           ,x"0008" -- 408E
           ,x"048a" -- 4090
           ,x"0028" -- 4092
           ,x"a3d8" -- 4094
           ,x"955e" -- 4096
           ,x"014e" -- 4098
           ,x"0220" -- 409A
           ,x"0028" -- 409C
           ,x"0028" -- 409E
           ,x"0024" -- 40A0
           ,x"9144" -- 40A2
           ,x"0028" -- 40A4
           ,x"036a" -- 40A6
           ,x"2d12" -- 40A8
           ,x"0160" -- 40AA
           ,x"0028" -- 40AC
           ,x"0028" -- 40AE
           ,x"0028" -- 40B0
           ,x"0020" -- 40B2
           ,x"0000" -- 40B4
           ,x"049e" -- 40B6
           ,x"0000" -- 40B8
           ,x"0000" -- 40BA
           ,x"0000" -- 40BC
           ,x"0000" -- 40BE
           ,x"0000" -- 40C0
           ,x"0000" -- 40C2
           ,x"0000" -- 40C4
           ,x"0000" -- 40C6
           ,x"0000" -- 40C8
           ,x"0000" -- 40CA
           ,x"0000" -- 40CC
           ,x"9882" -- 40CE
           ,x"9102" -- 40D0
           ,x"1cc2" -- 40D2
           ,x"7502" -- 40D4
           ,x"9bc6" -- 40D6
           ,x"860a" -- 40D8
           ,x"0c8c" -- 40DA
           ,x"a392" -- 40DC
           ,x"3bd8" -- 40DE
           ,x"c956" -- 40E0
           ,x"7266" -- 40E2
           ,x"9466" -- 40E4
           ,x"9e66" -- 40E6
           ,x"1a68" -- 40E8
           ,x"71e6" -- 40EA
           ,x"a244" -- 40EC
           ,x"1486" -- 40EE
           ,x"3486" -- 40F0
           ,x"695a" -- 40F2
           ,x"25da" -- 40F4
           ,x"7158" -- 40F6
           ,x"40da" -- 40F8
           ,x"9be0" -- 40FA
           ,x"63c6" -- 40FC
           ,x"23da" -- 40FE
           ,x"0000" -- 4100
           ,x"0000" -- 4102
           ,x"0000" -- 4104
           ,x"0000" -- 4106
           ,x"ffff" -- 4108
           ,x"4744" -- 410A
           ,x"3e43" -- 410C
           ,x"4248" -- 410E
           ,x"454c" -- 4110
           ,x"4d5f" -- 4112
           ,x"5d3f" -- 4114
           ,x"5c00" -- 4116
           ,x"5e00" -- 4118
           ,x"0000" -- 411A
           ,x"0000" -- 411C
           ,x"0000" -- 411E
           ,x"0000" -- 4120
           ,x"003c" -- 4122
           ,x"4059" -- 4124
           ,x"5657" -- 4126
           ,x"413d" -- 4128
           ,x"4c46" -- 412A
           ,x"4d60" -- 412C
           ,x"544f" -- 412E
           ,x"0038" -- 4130
           ,x"5441" -- 4132
           ,x"4200" -- 4134
           ,x"3953" -- 4136
           ,x"5445" -- 4138
           ,x"5000" -- 413A
           ,x"3a54" -- 413C
           ,x"4845" -- 413E
           ,x"4e00" -- 4140
           ,x"3b4f" -- 4142
           ,x"5200" -- 4144
           ,x"4e4c" -- 4146
           ,x"4f52" -- 4148
           ,x"004f" -- 414A
           ,x"414e" -- 414C
           ,x"4400" -- 414E
           ,x"504c" -- 4150
           ,x"414e" -- 4152
           ,x"4400" -- 4154
           ,x"514e" -- 4156
           ,x"4f54" -- 4158
           ,x"0052" -- 415A
           ,x"4c4e" -- 415C
           ,x"4f54" -- 415E
           ,x"0053" -- 4160
           ,x"4c58" -- 4162
           ,x"4f52" -- 4164
           ,x"0054" -- 4166
           ,x"003a" -- 4168
           ,x"4023" -- 416A
           ,x"2c3b" -- 416C
           ,x"3f25" -- 416E
           ,x"2422" -- 4170
           ,x"275c" -- 4172
           ,x"2126" -- 4174
           ,x"035b" -- 4176
           ,x"5d28" -- 4178
           ,x"291b" -- 417A
           ,x"6d4e" -- 417C
           ,x"6f38" -- 417E
           ,x"4208" -- 4180
           ,x"3d3d" -- 4182
           ,x"3e3e" -- 4184
           ,x"3c3c" -- 4186
           ,x"3c2d" -- 4188
           ,x"2b2f" -- 418A
           ,x"2a5e" -- 418C
           ,x"06a0" -- 418E
           ,x"a364" -- 4190
           ,x"0420" -- 4192
           ,x"8170" -- 4194
           ,x"04c1" -- 4196
           ,x"0706" -- 4198
           ,x"9838" -- 419A
           ,x"ab7f" -- 419C
           ,x"130e" -- 419E
           ,x"0608" -- 41A0
           ,x"06a0" -- 41A2
           ,x"b52a" -- 41A4
           ,x"1013" -- 41A6
           ,x"c820" -- 41A8
           ,x"801a" -- 41AA
           ,x"ef9e" -- 41AC
           ,x"0420" -- 41AE
           ,x"b558" -- 41B0
           ,x"0280" -- 41B2
           ,x"3800" -- 41B4
           ,x"1302" -- 41B6
           ,x"c181" -- 41B8
           ,x"1009" -- 41BA
           ,x"9838" -- 41BC
           ,x"c8bb" -- 41BE
           ,x"1306" -- 41C0
           ,x"0608" -- 41C2
           ,x"c820" -- 41C4
           ,x"8024" -- 41C6
           ,x"ef9e" -- 41C8
           ,x"0420" -- 41CA
           ,x"b558" -- 41CC
           ,x"c220" -- 41CE
           ,x"edd4" -- 41D0
           ,x"0648" -- 41D2
           ,x"8808" -- 41D4
           ,x"edd2" -- 41D6
           ,x"1217" -- 41D8
           ,x"0228" -- 41DA
           ,x"fffc" -- 41DC
           ,x"8601" -- 41DE
           ,x"15f9" -- 41E0
           ,x"0720" -- 41E2
           ,x"ede2" -- 41E4
           ,x"8808" -- 41E6
           ,x"edd2" -- 41E8
           ,x"1a0e" -- 41EA
           ,x"c078" -- 41EC
           ,x"8181" -- 41EE
           ,x"1b0b" -- 41F0
           ,x"06a0" -- 41F2
           ,x"ac2c" -- 41F4
           ,x"0420" -- 41F6
           ,x"8154" -- 41F8
           ,x"0228" -- 41FA
           ,x"fffa" -- 41FC
           ,x"0420" -- 41FE
           ,x"8190" -- 4200
           ,x"0420" -- 4202
           ,x"8170" -- 4204
           ,x"10ef" -- 4206
           ,x"0460" -- 4208
           ,x"8124" -- 420A
           ,x"dde0" -- 420C
           ,x"ab6c" -- 420E
           ,x"0583" -- 4210
           ,x"d073" -- 4212
           ,x"06c1" -- 4214
           ,x"d073" -- 4216
           ,x"06c1" -- 4218
           ,x"c820" -- 421A
           ,x"801a" -- 421C
           ,x"ef9e" -- 421E
           ,x"0420" -- 4220
           ,x"b05a" -- 4222
           ,x"9813" -- 4224
           ,x"c8c0" -- 4226
           ,x"13f1" -- 4228
           ,x"1055" -- 422A
           ,x"c28b" -- 422C
           ,x"0420" -- 422E
           ,x"81a4" -- 4230
           ,x"c1e0" -- 4232
           ,x"ed04" -- 4234
           ,x"c0d8" -- 4236
           ,x"a0e0" -- 4238
           ,x"ed0e" -- 423A
           ,x"020f" -- 423C
           ,x"2000" -- 423E
           ,x"ddcf" -- 4240
           ,x"c820" -- 4242
           ,x"801a" -- 4244
           ,x"ef9e" -- 4246
           ,x"0420" -- 4248
           ,x"b05a" -- 424A
           ,x"c0a0" -- 424C
           ,x"ede2" -- 424E
           ,x"9813" -- 4250
           ,x"ab76" -- 4252
           ,x"1601" -- 4254
           ,x"0642" -- 4256
           ,x"ddcf" -- 4258
           ,x"0582" -- 425A
           ,x"11fd" -- 425C
           ,x"9813" -- 425E
           ,x"ab81" -- 4260
           ,x"1601" -- 4262
           ,x"0607" -- 4264
           ,x"ddcf" -- 4266
           ,x"04c0" -- 4268
           ,x"d033" -- 426A
           ,x"0280" -- 426C
           ,x"0600" -- 426E
           ,x"131e" -- 4270
           ,x"0280" -- 4272
           ,x"4600" -- 4274
           ,x"1606" -- 4276
           ,x"dde0" -- 4278
           ,x"c8d6" -- 427A
           ,x"ddf3" -- 427C
           ,x"16fe" -- 427E
           ,x"0607" -- 4280
           ,x"100b" -- 4282
           ,x"0280" -- 4284
           ,x"4500" -- 4286
           ,x"1603" -- 4288
           ,x"dde0" -- 428A
           ,x"c8c0" -- 428C
           ,x"1005" -- 428E
           ,x"0280" -- 4290
           ,x"3f00" -- 4292
           ,x"1604" -- 4294
           ,x"dde0" -- 4296
           ,x"ab6d" -- 4298
           ,x"0870" -- 429A
           ,x"1003" -- 429C
           ,x"06a0" -- 429E
           ,x"ae62" -- 42A0
           ,x"a9b0" -- 42A2
           ,x"ddcf" -- 42A4
           ,x"0280" -- 42A6
           ,x"008e" -- 42A8
           ,x"1a01" -- 42AA
           ,x"0607" -- 42AC
           ,x"c380" -- 42AE
           ,x"0280" -- 42B0
           ,x"0006" -- 42B2
           ,x"11ae" -- 42B4
           ,x"13d8" -- 42B6
           ,x"0280" -- 42B8
           ,x"000a" -- 42BA
           ,x"1161" -- 42BC
           ,x"1502" -- 42BE
           ,x"0620" -- 42C0
           ,x"ede2" -- 42C2
           ,x"0280" -- 42C4
           ,x"0010" -- 42C6
           ,x"1605" -- 42C8
           ,x"05a0" -- 42CA
           ,x"ede2" -- 42CC
           ,x"1102" -- 42CE
           ,x"0720" -- 42D0
           ,x"ede2" -- 42D2
           ,x"c380" -- 42D4
           ,x"d033" -- 42D6
           ,x"133a" -- 42D8
           ,x"9800" -- 42DA
           ,x"c84e" -- 42DC
           ,x"1a5d" -- 42DE
           ,x"9800" -- 42E0
           ,x"ab7f" -- 42E2
           ,x"1a61" -- 42E4
           ,x"0980" -- 42E6
           ,x"c100" -- 42E8
           ,x"0280" -- 42EA
           ,x"003c" -- 42EC
           ,x"1a66" -- 42EE
           ,x"0280" -- 42F0
           ,x"004e" -- 42F2
           ,x"1a03" -- 42F4
           ,x"0280" -- 42F6
           ,x"0054" -- 42F8
           ,x"125e" -- 42FA
           ,x"0280" -- 42FC
           ,x"0062" -- 42FE
           ,x"1a28" -- 4300
           ,x"0280" -- 4302
           ,x"006f" -- 4304
           ,x"1a65" -- 4306
           ,x"137b" -- 4308
           ,x"c160" -- 430A
           ,x"edd4" -- 430C
           ,x"a000" -- 430E
           ,x"a140" -- 4310
           ,x"04c2" -- 4312
           ,x"c165" -- 4314
           ,x"ff20" -- 4316
           ,x"1503" -- 4318
           ,x"0505" -- 431A
           ,x"0202" -- 431C
           ,x"004a" -- 431E
           ,x"2160" -- 4320
           ,x"a56e" -- 4322
           ,x"160c" -- 4324
           ,x"06a0" -- 4326
           ,x"ae88" -- 4328
           ,x"0921" -- 432A
           ,x"c045" -- 432C
           ,x"0241" -- 432E
           ,x"007f" -- 4330
           ,x"c820" -- 4332
           ,x"801a" -- 4334
           ,x"ef9e" -- 4336
           ,x"0420" -- 4338
           ,x"b05a" -- 433A
           ,x"1005" -- 433C
           ,x"0a15" -- 433E
           ,x"020d" -- 4340
           ,x"ad48" -- 4342
           ,x"0460" -- 4344
           ,x"ae6c" -- 4346
           ,x"c102" -- 4348
           ,x"162b" -- 434A
           ,x"10c4" -- 434C
           ,x"75d7" -- 434E
           ,x"045a" -- 4350
           ,x"dde4" -- 4352
           ,x"ab2d" -- 4354
           ,x"06c0" -- 4356
           ,x"06a0" -- 4358
           ,x"872c" -- 435A
           ,x"2044" -- 435C
           ,x"2045" -- 435E
           ,x"0c47" -- 4360
           ,x"1d3c" -- 4362
           ,x"0000" -- 4364
           ,x"06a0" -- 4366
           ,x"ad8a" -- 4368
           ,x"3d55" -- 436A
           ,x"3d58" -- 436C
           ,x"3d5a" -- 436E
           ,x"3e5b" -- 4370
           ,x"0000" -- 4372
           ,x"0607" -- 4374
           ,x"ddcf" -- 4376
           ,x"ddcf" -- 4378
           ,x"dde4" -- 437A
           ,x"ab2d" -- 437C
           ,x"1001" -- 437E
           ,x"0607" -- 4380
           ,x"ddf3" -- 4382
           ,x"16fe" -- 4384
           ,x"0607" -- 4386
           ,x"045a" -- 4388
           ,x"d5fb" -- 438A
           ,x"13a4" -- 438C
           ,x"9ec0" -- 438E
           ,x"16fc" -- 4390
           ,x"0587" -- 4392
           ,x"10a0" -- 4394
           ,x"0460" -- 4396
           ,x"ac66" -- 4398
           ,x"1039" -- 439A
           ,x"ddf3" -- 439C
           ,x"16fe" -- 439E
           ,x"0607" -- 43A0
           ,x"dde4" -- 43A2
           ,x"ab2d" -- 43A4
           ,x"1097" -- 43A6
           ,x"06a0" -- 43A8
           ,x"ae62" -- 43AA
           ,x"aa98" -- 43AC
           ,x"9813" -- 43AE
           ,x"ad1f" -- 43B0
           ,x"1391" -- 43B2
           ,x"ddcf" -- 43B4
           ,x"108f" -- 43B6
           ,x"0224" -- 43B8
           ,x"ffee" -- 43BA
           ,x"ddcf" -- 43BC
           ,x"a104" -- 43BE
           ,x"c164" -- 43C0
           ,x"addc" -- 43C2
           ,x"ddf5" -- 43C4
           ,x"d015" -- 43C6
           ,x"16fd" -- 43C8
           ,x"0284" -- 43CA
           ,x"0076" -- 43CC
           ,x"13e3" -- 43CE
           ,x"10f1" -- 43D0
           ,x"0280" -- 43D2
           ,x"006d" -- 43D4
           ,x"1404" -- 43D6
           ,x"0220" -- 43D8
           ,x"ff9d" -- 43DA
           ,x"c040" -- 43DC
           ,x"1007" -- 43DE
           ,x"d073" -- 43E0
           ,x"06c1" -- 43E2
           ,x"d073" -- 43E4
           ,x"06c1" -- 43E6
           ,x"0280" -- 43E8
           ,x"006e" -- 43EA
           ,x"1306" -- 43EC
           ,x"c820" -- 43EE
           ,x"801a" -- 43F0
           ,x"ef9e" -- 43F2
           ,x"0420" -- 43F4
           ,x"b05a" -- 43F6
           ,x"10de" -- 43F8
           ,x"06a0" -- 43FA
           ,x"9c8e" -- 43FC
           ,x"10db" -- 43FE
           ,x"c803" -- 4400
           ,x"ef9e" -- 4402
           ,x"0420" -- 4404
           ,x"b05e" -- 4406
           ,x"0223" -- 4408
           ,x"0006" -- 440A
           ,x"10d4" -- 440C
           ,x"dde0" -- 440E
           ,x"ab2b" -- 4410
           ,x"dde0" -- 4412
           ,x"ab7d" -- 4414
           ,x"0220" -- 4416
           ,x"4000" -- 4418
           ,x"ddc0" -- 441A
           ,x"028e" -- 441C
           ,x"0084" -- 441E
           ,x"16c6" -- 4420
           ,x"c3a0" -- 4422
           ,x"edd4" -- 4424
           ,x"9813" -- 4426
           ,x"ab26" -- 4428
           ,x"13c5" -- 442A
           ,x"dde0" -- 442C
           ,x"ab77" -- 442E
           ,x"d7b3" -- 4430
           ,x"c07e" -- 4432
           ,x"0821" -- 4434
           ,x"06a0" -- 4436
           ,x"ae92" -- 4438
           ,x"9813" -- 443A
           ,x"ab26" -- 443C
           ,x"1303" -- 443E
           ,x"dde0" -- 4440
           ,x"ab6c" -- 4442
           ,x"10f5" -- 4444
           ,x"dde0" -- 4446
           ,x"ab78" -- 4448
           ,x"10b5" -- 444A
           ,x"ab2e" -- 444C
           ,x"ab32" -- 444E
           ,x"ab37" -- 4450
           ,x"ab3d" -- 4452
           ,x"ab43" -- 4454
           ,x"ab47" -- 4456
           ,x"ab4c" -- 4458
           ,x"ab51" -- 445A
           ,x"ab57" -- 445C
           ,x"ab5c" -- 445E
           ,x"ab62" -- 4460
           ,x"c13b" -- 4462
           ,x"c34b" -- 4464
           ,x"0870" -- 4466
           ,x"a100" -- 4468
           ,x"c154" -- 446A
           ,x"06a0" -- 446C
           ,x"ae88" -- 446E
           ,x"0a71" -- 4470
           ,x"06a0" -- 4472
           ,x"ae88" -- 4474
           ,x"0a21" -- 4476
           ,x"06a0" -- 4478
           ,x"ae88" -- 447A
           ,x"0931" -- 447C
           ,x"0224" -- 447E
           ,x"00ac" -- 4480
           ,x"0915" -- 4482
           ,x"18f2" -- 4484
           ,x"045d" -- 4486
           ,x"c045" -- 4488
           ,x"04bb" -- 448A
           ,x"0241" -- 448C
           ,x"1f00" -- 448E
           ,x"1303" -- 4490
           ,x"0221" -- 4492
           ,x"4000" -- 4494
           ,x"ddc1" -- 4496
           ,x"045b" -- 4498
           ,x"c820" -- 449A
           ,x"ed04" -- 449C
           ,x"edda" -- 449E
           ,x"c820" -- 44A0
           ,x"ed0a" -- 44A2
           ,x"eddc" -- 44A4
           ,x"04f1" -- 44A6
           ,x"0281" -- 44A8
           ,x"ed00" -- 44AA
           ,x"1afc" -- 44AC
           ,x"04e0" -- 44AE
           ,x"ed2a" -- 44B0
           ,x"c820" -- 44B2
           ,x"edd4" -- 44B4
           ,x"edea" -- 44B6
           ,x"04e0" -- 44B8
           ,x"edec" -- 44BA
           ,x"045b" -- 44BC
           ,x"0420" -- 44BE
           ,x"8170" -- 44C0
           ,x"0720" -- 44C2
           ,x"ede4" -- 44C4
           ,x"04e0" -- 44C6
           ,x"8046" -- 44C8
           ,x"c820" -- 44CA
           ,x"edd4" -- 44CC
           ,x"ede6" -- 44CE
           ,x"c060" -- 44D0
           ,x"edd6" -- 44D2
           ,x"06a0" -- 44D4
           ,x"ae9a" -- 44D6
           ,x"1014" -- 44D8
           ,x"0280" -- 44DA
           ,x"3c00" -- 44DC
           ,x"1603" -- 44DE
           ,x"05a0" -- 44E0
           ,x"ed12" -- 44E2
           ,x"1029" -- 44E4
           ,x"0280" -- 44E6
           ,x"3b00" -- 44E8
           ,x"1326" -- 44EA
           ,x"0280" -- 44EC
           ,x"4700" -- 44EE
           ,x"1308" -- 44F0
           ,x"0420" -- 44F2
           ,x"8d70" -- 44F4
           ,x"0025" -- 44F6
           ,x"d838" -- 44F8
           ,x"ede8" -- 44FA
           ,x"c020" -- 44FC
           ,x"ede8" -- 44FE
           ,x"16ec" -- 4500
           ,x"c220" -- 4502
           ,x"8046" -- 4504
           ,x"1607" -- 4506
           ,x"0420" -- 4508
           ,x"8194" -- 450A
           ,x"1000" -- 450C
           ,x"1000" -- 450E
           ,x"c020" -- 4510
           ,x"ede4" -- 4512
           ,x"134a" -- 4514
           ,x"c220" -- 4516
           ,x"ede6" -- 4518
           ,x"0228" -- 451A
           ,x"fffc" -- 451C
           ,x"8808" -- 451E
           ,x"edd2" -- 4520
           ,x"1a45" -- 4522
           ,x"c808" -- 4524
           ,x"ede6" -- 4526
           ,x"c828" -- 4528
           ,x"fffe" -- 452A
           ,x"ed32" -- 452C
           ,x"c218" -- 452E
           ,x"a220" -- 4530
           ,x"ed0e" -- 4532
           ,x"04e0" -- 4534
           ,x"ed12" -- 4536
           ,x"04e0" -- 4538
           ,x"edf0" -- 453A
           ,x"04c2" -- 453C
           ,x"d0b8" -- 453E
           ,x"0972" -- 4540
           ,x"0282" -- 4542
           ,x"0096" -- 4544
           ,x"1b2e" -- 4546
           ,x"c262" -- 4548
           ,x"afba" -- 454A
           ,x"132b" -- 454C
           ,x"c2e0" -- 454E
           ,x"ed30" -- 4550
           ,x"1327" -- 4552
           ,x"c2e0" -- 4554
           ,x"ede4" -- 4556
           ,x"1324" -- 4558
           ,x"06a0" -- 455A
           ,x"a214" -- 455C
           ,x"2053" -- 455E
           ,x"7461" -- 4560
           ,x"7465" -- 4562
           ,x"6d65" -- 4564
           ,x"6e74" -- 4566
           ,x"204e" -- 4568
           ,x"6f2e" -- 456A
           ,x"2000" -- 456C
           ,x"c2e0" -- 456E
           ,x"ede6" -- 4570
           ,x"c80b" -- 4572
           ,x"ef9e" -- 4574
           ,x"0660" -- 4576
           ,x"ef9e" -- 4578
           ,x"0420" -- 457A
           ,x"b05a" -- 457C
           ,x"c2e0" -- 457E
           ,x"ed12" -- 4580
           ,x"1307" -- 4582
           ,x"dde0" -- 4584
           ,x"c875" -- 4586
           ,x"c820" -- 4588
           ,x"8026" -- 458A
           ,x"ef9e" -- 458C
           ,x"0420" -- 458E
           ,x"b05a" -- 4590
           ,x"06a0" -- 4592
           ,x"a218" -- 4594
           ,x"2020" -- 4596
           ,x"2000" -- 4598
           ,x"0420" -- 459A
           ,x"8190" -- 459C
           ,x"0420" -- 459E
           ,x"8170" -- 45A0
           ,x"0459" -- 45A2
           ,x"0420" -- 45A4
           ,x"8d70" -- 45A6
           ,x"ffff" -- 45A8
           ,x"0460" -- 45AA
           ,x"8124" -- 45AC
           ,x"0460" -- 45AE
           ,x"8dde" -- 45B0
           ,x"c020" -- 45B2
           ,x"ed38" -- 45B4
           ,x"16c0" -- 45B6
           ,x"10a4" -- 45B8
           ,x"8dde" -- 45BA
           ,x"950e" -- 45BC
           ,x"9512" -- 45BE
           ,x"afb2" -- 45C0
           ,x"af02" -- 45C2
           ,x"9100" -- 45C4
           ,x"97b8" -- 45C6
           ,x"af02" -- 45C8
           ,x"9206" -- 45CA
           ,x"8e38" -- 45CC
           ,x"9b6e" -- 45CE
           ,x"8ebc" -- 45D0
           ,x"8748" -- 45D2
           ,x"9654" -- 45D4
           ,x"9df4" -- 45D6
           ,x"9e30" -- 45D8
           ,x"9588" -- 45DA
           ,x"8dc4" -- 45DC
           ,x"a260" -- 45DE
           ,x"a24c" -- 45E0
           ,x"8742" -- 45E2
           ,x"8f38" -- 45E4
           ,x"90f2" -- 45E6
           ,x"90f8" -- 45E8
           ,x"9d88" -- 45EA
           ,x"80b6" -- 45EC
           ,x"90ae" -- 45EE
           ,x"c334" -- 45F0
           ,x"c330" -- 45F2
           ,x"8a38" -- 45F4
           ,x"9cd4" -- 45F6
           ,x"89dc" -- 45F8
           ,x"89d4" -- 45FA
           ,x"8ac6" -- 45FC
           ,x"89e2" -- 45FE
           ,x"9a50" -- 4600
           ,x"ab8e" -- 4602
           ,x"9e7a" -- 4604
           ,x"8b28" -- 4606
           ,x"8ae0" -- 4608
           ,x"8946" -- 460A
           ,x"88cc" -- 460C
           ,x"a2a0" -- 460E
           ,x"a2be" -- 4610
           ,x"0000" -- 4612
           ,x"874e" -- 4614
           ,x"0000" -- 4616
           ,x"0000" -- 4618
           ,x"0000" -- 461A
           ,x"0000" -- 461C
           ,x"0000" -- 461E
           ,x"0000" -- 4620
           ,x"0000" -- 4622
           ,x"0000" -- 4624
           ,x"0000" -- 4626
           ,x"0000" -- 4628
           ,x"0000" -- 462A
           ,x"8ba8" -- 462C
           ,x"a25a" -- 462E
           ,x"a252" -- 4630
           ,x"95b8" -- 4632
           ,x"8fe4" -- 4634
           ,x"97b8" -- 4636
           ,x"9b6e" -- 4638
           ,x"9a8c" -- 463A
           ,x"95ca" -- 463C
           ,x"8fc0" -- 463E
           ,x"80c4" -- 4640
           ,x"8dde" -- 4642
           ,x"9b6e" -- 4644
           ,x"c72e" -- 4646
           ,x"bfa8" -- 4648
           ,x"8f5e" -- 464A
           ,x"8f44" -- 464C
           ,x"9984" -- 464E
           ,x"9a1e" -- 4650
           ,x"0700" -- 4652
           ,x"0420" -- 4654
           ,x"8d70" -- 4656
           ,x"0022" -- 4658
           ,x"ef88" -- 465A
           ,x"b062" -- 465C
           ,x"ef88" -- 465E
           ,x"b06c" -- 4660
           ,x"0420" -- 4662
           ,x"be74" -- 4664
           ,x"c81b" -- 4666
           ,x"ef6a" -- 4668
           ,x"1008" -- 466A
           ,x"020a" -- 466C
           ,x"ef68" -- 466E
           ,x"debb" -- 4670
           ,x"debb" -- 4672
           ,x"debb" -- 4674
           ,x"debb" -- 4676
           ,x"debb" -- 4678
           ,x"d69b" -- 467A
           ,x"0420" -- 467C
           ,x"bd1a" -- 467E
           ,x"04cc" -- 4680
           ,x"0207" -- 4682
           ,x"edfe" -- 4684
           ,x"7dd7" -- 4686
           ,x"c060" -- 4688
           ,x"ef68" -- 468A
           ,x"1106" -- 468C
           ,x"1508" -- 468E
           ,x"dde0" -- 4690
           ,x"b0f7" -- 4692
           ,x"020a" -- 4694
           ,x"000c" -- 4696
           ,x"1046" -- 4698
           ,x"0420" -- 469A
           ,x"bd0c" -- 469C
           ,x"070c" -- 469E
           ,x"0241" -- 46A0
           ,x"00f0" -- 46A2
           ,x"13d7" -- 46A4
           ,x"04ca" -- 46A6
           ,x"d060" -- 46A8
           ,x"ef68" -- 46AA
           ,x"0981" -- 46AC
           ,x"0208" -- 46AE
           ,x"004a" -- 46B0
           ,x"6201" -- 46B2
           ,x"1316" -- 46B4
           ,x"1108" -- 46B6
           ,x"06a0" -- 46B8
           ,x"b48a" -- 46BA
           ,x"a288" -- 46BC
           ,x"c800" -- 46BE
           ,x"ef7e" -- 46C0
           ,x"0420" -- 46C2
           ,x"bd84" -- 46C4
           ,x"10f0" -- 46C6
           ,x"0508" -- 46C8
           ,x"06a0" -- 46CA
           ,x"b48a" -- 46CC
           ,x"6288" -- 46CE
           ,x"c800" -- 46D0
           ,x"ef7e" -- 46D2
           ,x"0420" -- 46D4
           ,x"beac" -- 46D6
           ,x"10e7" -- 46D8
           ,x"06a0" -- 46DA
           ,x"bf54" -- 46DC
           ,x"058a" -- 46DE
           ,x"100b" -- 46E0
           ,x"c820" -- 46E2
           ,x"8016" -- 46E4
           ,x"ef7e" -- 46E6
           ,x"0420" -- 46E8
           ,x"bc32" -- 46EA
           ,x"0240" -- 46EC
           ,x"00ff" -- 46EE
           ,x"0203" -- 46F0
           ,x"b236" -- 46F2
           ,x"0209" -- 46F4
           ,x"0030" -- 46F6
           ,x"c133" -- 46F8
           ,x"c173" -- 46FA
           ,x"c1b3" -- 46FC
           ,x"06a0" -- 46FE
           ,x"bf68" -- 4700
           ,x"11eb" -- 4702
           ,x"0589" -- 4704
           ,x"06a0" -- 4706
           ,x"bf68" -- 4708
           ,x"13fc" -- 470A
           ,x"15fb" -- 470C
           ,x"06a0" -- 470E
           ,x"bf54" -- 4710
           ,x"06c9" -- 4712
           ,x"ddc9" -- 4714
           ,x"0209" -- 4716
           ,x"002f" -- 4718
           ,x"c133" -- 471A
           ,x"c173" -- 471C
           ,x"c1b3" -- 471E
           ,x"0283" -- 4720
           ,x"b284" -- 4722
           ,x"12ef" -- 4724
           ,x"7dd7" -- 4726
           ,x"0287" -- 4728
           ,x"ee0d" -- 472A
           ,x"1afc" -- 472C
           ,x"c1ed" -- 472E
           ,x"000e" -- 4730
           ,x"0200" -- 4732
           ,x"000a" -- 4734
           ,x"c260" -- 4736
           ,x"ed3a" -- 4738
           ,x"160a" -- 473A
           ,x"06a0" -- 473C
           ,x"b1e8" -- 473E
           ,x"060a" -- 4740
           ,x"04c4" -- 4742
           ,x"9560" -- 4744
           ,x"b0f7" -- 4746
           ,x"1605" -- 4748
           ,x"d544" -- 474A
           ,x"0605" -- 474C
           ,x"10fa" -- 474E
           ,x"0460" -- 4750
           ,x"92a8" -- 4752
           ,x"c30c" -- 4754
           ,x"1302" -- 4756
           ,x"dde0" -- 4758
           ,x"c8c7" -- 475A
           ,x"064a" -- 475C
           ,x"1127" -- 475E
           ,x"028a" -- 4760
           ,x"0010" -- 4762
           ,x"1524" -- 4764
           ,x"022a" -- 4766
           ,x"fff5" -- 4768
           ,x"1510" -- 476A
           ,x"130f" -- 476C
           ,x"ddf3" -- 476E
           ,x"1307" -- 4770
           ,x"058a" -- 4772
           ,x"11fc" -- 4774
           ,x"d013" -- 4776
           ,x"1315" -- 4778
           ,x"dde0" -- 477A
           ,x"c875" -- 477C
           ,x"100f" -- 477E
           ,x"0607" -- 4780
           ,x"dde0" -- 4782
           ,x"b0f7" -- 4784
           ,x"058a" -- 4786
           ,x"11fc" -- 4788
           ,x"100c" -- 478A
           ,x"dde0" -- 478C
           ,x"b0f7" -- 478E
           ,x"dde0" -- 4790
           ,x"c875" -- 4792
           ,x"060a" -- 4794
           ,x"1103" -- 4796
           ,x"dde0" -- 4798
           ,x"b0f7" -- 479A
           ,x"10fb" -- 479C
           ,x"ddf3" -- 479E
           ,x"16fe" -- 47A0
           ,x"0607" -- 47A2
           ,x"cb47" -- 47A4
           ,x"000e" -- 47A6
           ,x"0380" -- 47A8
           ,x"c1c6" -- 47AA
           ,x"10fb" -- 47AC
           ,x"ddf3" -- 47AE
           ,x"d113" -- 47B0
           ,x"1302" -- 47B2
           ,x"dde0" -- 47B4
           ,x"c875" -- 47B6
           ,x"ddf3" -- 47B8
           ,x"16fe" -- 47BA
           ,x"0607" -- 47BC
           ,x"dde0" -- 47BE
           ,x"c842" -- 47C0
           ,x"022a" -- 47C2
           ,x"fff6" -- 47C4
           ,x"050a" -- 47C6
           ,x"1503" -- 47C8
           ,x"dde0" -- 47CA
           ,x"c8c7" -- 47CC
           ,x"050a" -- 47CE
           ,x"04c9" -- 47D0
           ,x"3e60" -- 47D2
           ,x"b27c" -- 47D4
           ,x"0229" -- 47D6
           ,x"0030" -- 47D8
           ,x"022a" -- 47DA
           ,x"0030" -- 47DC
           ,x"06c9" -- 47DE
           ,x"06ca" -- 47E0
           ,x"ddc9" -- 47E2
           ,x"ddca" -- 47E4
           ,x"10de" -- 47E6
           ,x"0206" -- 47E8
           ,x"edff" -- 47EA
           ,x"d820" -- 47EC
           ,x"b0f7" -- 47EE
           ,x"ee0a" -- 47F0
           ,x"a180" -- 47F2
           ,x"d000" -- 47F4
           ,x"1618" -- 47F6
           ,x"c146" -- 47F8
           ,x"0586" -- 47FA
           ,x"d0d6" -- 47FC
           ,x"1314" -- 47FE
           ,x"d580" -- 4800
           ,x"b0e0" -- 4802
           ,x"b925" -- 4804
           ,x"90e0" -- 4806
           ,x"c8dd" -- 4808
           ,x"1b0e" -- 480A
           ,x"0606" -- 480C
           ,x"d016" -- 480E
           ,x"1308" -- 4810
           ,x"b5a0" -- 4812
           ,x"b921" -- 4814
           ,x"95a0" -- 4816
           ,x"c8dd" -- 4818
           ,x"1b06" -- 481A
           ,x"d5a0" -- 481C
           ,x"b0f7" -- 481E
           ,x"10f5" -- 4820
           ,x"049b" -- 4822
           ,x"d5a0" -- 4824
           ,x"c84d" -- 4826
           ,x"0203" -- 4828
           ,x"edfe" -- 482A
           ,x"d1b3" -- 482C
           ,x"1301" -- 482E
           ,x"0603" -- 4830
           ,x"046b" -- 4832
           ,x"0002" -- 4834
           ,x"00e8" -- 4836
           ,x"d4a5" -- 4838
           ,x"1000" -- 483A
           ,x"0017" -- 483C
           ,x"4876" -- 483E
           ,x"e800" -- 4840
           ,x"0002" -- 4842
           ,x"540b" -- 4844
           ,x"e400" -- 4846
           ,x"0000" -- 4848
           ,x"3b9a" -- 484A
           ,x"ca00" -- 484C
           ,x"0000" -- 484E
           ,x"05f5" -- 4850
           ,x"e100" -- 4852
           ,x"0000" -- 4854
           ,x"0098" -- 4856
           ,x"9680" -- 4858
           ,x"0000" -- 485A
           ,x"000f" -- 485C
           ,x"4240" -- 485E
           ,x"0000" -- 4860
           ,x"0001" -- 4862
           ,x"86a0" -- 4864
           ,x"0000" -- 4866
           ,x"0000" -- 4868
           ,x"2710" -- 486A
           ,x"0000" -- 486C
           ,x"0000" -- 486E
           ,x"03e8" -- 4870
           ,x"0000" -- 4872
           ,x"0000" -- 4874
           ,x"0064" -- 4876
           ,x"0000" -- 4878
           ,x"0000" -- 487A
           ,x"000a" -- 487C
           ,x"0000" -- 487E
           ,x"0000" -- 4880
           ,x"0001" -- 4882
           ,x"ef88" -- 4884
           ,x"b28c" -- 4886
           ,x"ef88" -- 4888
           ,x"b290" -- 488A
           ,x"04c8" -- 488C
           ,x"1001" -- 488E
           ,x"0708" -- 4890
           ,x"c1ed" -- 4892
           ,x"000e" -- 4894
           ,x"04c2" -- 4896
           ,x"04c4" -- 4898
           ,x"06a0" -- 489A
           ,x"b436" -- 489C
           ,x"103a" -- 489E
           ,x"0704" -- 48A0
           ,x"c187" -- 48A2
           ,x"d036" -- 48A4
           ,x"0980" -- 48A6
           ,x"0220" -- 48A8
           ,x"ffd0" -- 48AA
           ,x"1114" -- 48AC
           ,x"0280" -- 48AE
           ,x"0009" -- 48B0
           ,x"1208" -- 48B2
           ,x"0220" -- 48B4
           ,x"fff9" -- 48B6
           ,x"0280" -- 48B8
           ,x"000a" -- 48BA
           ,x"110c" -- 48BC
           ,x"0280" -- 48BE
           ,x"000f" -- 48C0
           ,x"1b03" -- 48C2
           ,x"0a42" -- 48C4
           ,x"a080" -- 48C6
           ,x"10ed" -- 48C8
           ,x"0220" -- 48CA
           ,x"ffef" -- 48CC
           ,x"1603" -- 48CE
           ,x"d036" -- 48D0
           ,x"c1c6" -- 48D2
           ,x"1017" -- 48D4
           ,x"04c2" -- 48D6
           ,x"06a0" -- 48D8
           ,x"b416" -- 48DA
           ,x"100a" -- 48DC
           ,x"c042" -- 48DE
           ,x"3860" -- 48E0
           ,x"b27c" -- 48E2
           ,x"c041" -- 48E4
           ,x"161b" -- 48E6
           ,x"c082" -- 48E8
           ,x"1119" -- 48EA
           ,x"a080" -- 48EC
           ,x"1117" -- 48EE
           ,x"10f3" -- 48F0
           ,x"0280" -- 48F2
           ,x"2e00" -- 48F4
           ,x"1311" -- 48F6
           ,x"0280" -- 48F8
           ,x"4500" -- 48FA
           ,x"130e" -- 48FC
           ,x"c208" -- 48FE
           ,x"1301" -- 4900
           ,x"05ce" -- 4902
           ,x"c104" -- 4904
           ,x"1301" -- 4906
           ,x"0502" -- 4908
           ,x"cb42" -- 490A
           ,x"0002" -- 490C
           ,x"cb47" -- 490E
           ,x"000e" -- 4910
           ,x"05ce" -- 4912
           ,x"05ce" -- 4914
           ,x"c740" -- 4916
           ,x"0380" -- 4918
           ,x"c208" -- 491A
           ,x"13f3" -- 491C
           ,x"0420" -- 491E
           ,x"be74" -- 4920
           ,x"c1ed" -- 4922
           ,x"000e" -- 4924
           ,x"0702" -- 4926
           ,x"04c6" -- 4928
           ,x"04cc" -- 492A
           ,x"04c4" -- 492C
           ,x"06a0" -- 492E
           ,x"b436" -- 4930
           ,x"10f0" -- 4932
           ,x"070c" -- 4934
           ,x"06a0" -- 4936
           ,x"b416" -- 4938
           ,x"101d" -- 493A
           ,x"c082" -- 493C
           ,x"1101" -- 493E
           ,x"0586" -- 4940
           ,x"c000" -- 4942
           ,x"1602" -- 4944
           ,x"c104" -- 4946
           ,x"13f6" -- 4948
           ,x"0584" -- 494A
           ,x"0284" -- 494C
           ,x"000b" -- 494E
           ,x"1201" -- 4950
           ,x"04c0" -- 4952
           ,x"c820" -- 4954
           ,x"800c" -- 4956
           ,x"ef7e" -- 4958
           ,x"0420" -- 495A
           ,x"bd84" -- 495C
           ,x"0a40" -- 495E
           ,x"13ea" -- 4960
           ,x"0220" -- 4962
           ,x"4100" -- 4964
           ,x"c800" -- 4966
           ,x"edf8" -- 4968
           ,x"c820" -- 496A
           ,x"800a" -- 496C
           ,x"ef7e" -- 496E
           ,x"0420" -- 4970
           ,x"bc4a" -- 4972
           ,x"10e0" -- 4974
           ,x"0280" -- 4976
           ,x"2e00" -- 4978
           ,x"1606" -- 497A
           ,x"c082" -- 497C
           ,x"1319" -- 497E
           ,x"c208" -- 4980
           ,x"1317" -- 4982
           ,x"04c2" -- 4984
           ,x"10d7" -- 4986
           ,x"0280" -- 4988
           ,x"4500" -- 498A
           ,x"1612" -- 498C
           ,x"0205" -- 498E
           ,x"0501" -- 4990
           ,x"06a0" -- 4992
           ,x"b436" -- 4994
           ,x"10be" -- 4996
           ,x"0ac5" -- 4998
           ,x"04c1" -- 499A
           ,x"06a0" -- 499C
           ,x"b416" -- 499E
           ,x"1006" -- 49A0
           ,x"c0c1" -- 49A2
           ,x"38e0" -- 49A4
           ,x"b27c" -- 49A6
           ,x"a100" -- 49A8
           ,x"c044" -- 49AA
           ,x"10f7" -- 49AC
           ,x"0485" -- 49AE
           ,x"a181" -- 49B0
           ,x"c740" -- 49B2
           ,x"cb47" -- 49B4
           ,x"000e" -- 49B6
           ,x"c206" -- 49B8
           ,x"1109" -- 49BA
           ,x"1311" -- 49BC
           ,x"06a0" -- 49BE
           ,x"b492" -- 49C0
           ,x"6188" -- 49C2
           ,x"c800" -- 49C4
           ,x"ef7e" -- 49C6
           ,x"0420" -- 49C8
           ,x"beac" -- 49CA
           ,x"10f5" -- 49CC
           ,x"0508" -- 49CE
           ,x"06a0" -- 49D0
           ,x"b492" -- 49D2
           ,x"a188" -- 49D4
           ,x"c800" -- 49D6
           ,x"ef7e" -- 49D8
           ,x"0420" -- 49DA
           ,x"bd84" -- 49DC
           ,x"10ec" -- 49DE
           ,x"c30c" -- 49E0
           ,x"1314" -- 49E2
           ,x"0420" -- 49E4
           ,x"bd0c" -- 49E6
           ,x"020c" -- 49E8
           ,x"ef68" -- 49EA
           ,x"c0cc" -- 49EC
           ,x"0206" -- 49EE
           ,x"b40e" -- 49F0
           ,x"8dbc" -- 49F2
           ,x"160b" -- 49F4
           ,x"8dbc" -- 49F6
           ,x"1609" -- 49F8
           ,x"8d9c" -- 49FA
           ,x"1607" -- 49FC
           ,x"04f3" -- 49FE
           ,x"ccd6" -- 4A00
           ,x"c096" -- 4A02
           ,x"04d3" -- 4A04
           ,x"04c4" -- 4A06
           ,x"0460" -- 4A08
           ,x"b2fe" -- 4A0A
           ,x"0380" -- 4A0C
           ,x"c480" -- 4A0E
           ,x"0000" -- 4A10
           ,x"0000" -- 4A12
           ,x"8000" -- 4A14
           ,x"04c0" -- 4A16
           ,x"d037" -- 4A18
           ,x"130c" -- 4A1A
           ,x"0280" -- 4A1C
           ,x"2000" -- 4A1E
           ,x"13fa" -- 4A20
           ,x"0280" -- 4A22
           ,x"3000" -- 4A24
           ,x"1a06" -- 4A26
           ,x"0280" -- 4A28
           ,x"3900" -- 4A2A
           ,x"1b03" -- 4A2C
           ,x"0a40" -- 4A2E
           ,x"09c0" -- 4A30
           ,x"05cb" -- 4A32
           ,x"045b" -- 4A34
           ,x"9837" -- 4A36
           ,x"c0e4" -- 4A38
           ,x"13fd" -- 4A3A
           ,x"0607" -- 4A3C
           ,x"c047" -- 4A3E
           ,x"c28b" -- 4A40
           ,x"06a0" -- 4A42
           ,x"b416" -- 4A44
           ,x"1004" -- 4A46
           ,x"05ca" -- 4A48
           ,x"05ca" -- 4A4A
           ,x"c1c1" -- 4A4C
           ,x"045a" -- 4A4E
           ,x"0280" -- 4A50
           ,x"2b00" -- 4A52
           ,x"1307" -- 4A54
           ,x"0280" -- 4A56
           ,x"2d00" -- 4A58
           ,x"1307" -- 4A5A
           ,x"0280" -- 4A5C
           ,x"2e00" -- 4A5E
           ,x"16f5" -- 4A60
           ,x"0607" -- 4A62
           ,x"06a0" -- 4A64
           ,x"b470" -- 4A66
           ,x"10ef" -- 4A68
           ,x"06a0" -- 4A6A
           ,x"b470" -- 4A6C
           ,x"10ed" -- 4A6E
           ,x"c0cb" -- 4A70
           ,x"c047" -- 4A72
           ,x"06a0" -- 4A74
           ,x"b416" -- 4A76
           ,x"1001" -- 4A78
           ,x"0453" -- 4A7A
           ,x"0280" -- 4A7C
           ,x"2e00" -- 4A7E
           ,x"16e5" -- 4A80
           ,x"06a0" -- 4A82
           ,x"b416" -- 4A84
           ,x"10e2" -- 4A86
           ,x"0453" -- 4A88
           ,x"0288" -- 4A8A
           ,x"0005" -- 4A8C
           ,x"1a06" -- 4A8E
           ,x"0588" -- 4A90
           ,x"0288" -- 4A92
           ,x"000a" -- 4A94
           ,x"1a02" -- 4A96
           ,x"0208" -- 4A98
           ,x"0009" -- 4A9A
           ,x"04bb" -- 4A9C
           ,x"0200" -- 4A9E
           ,x"b4ac" -- 4AA0
           ,x"0a18" -- 4AA2
           ,x"a008" -- 4AA4
           ,x"0a18" -- 4AA6
           ,x"a008" -- 4AA8
           ,x"045b" -- 4AAA
           ,x"4110" -- 4AAC
           ,x"0000" -- 4AAE
           ,x"0000" -- 4AB0
           ,x"41a0" -- 4AB2
           ,x"0000" -- 4AB4
           ,x"0000" -- 4AB6
           ,x"4264" -- 4AB8
           ,x"0000" -- 4ABA
           ,x"0000" -- 4ABC
           ,x"433e" -- 4ABE
           ,x"8000" -- 4AC0
           ,x"0000" -- 4AC2
           ,x"4427" -- 4AC4
           ,x"1000" -- 4AC6
           ,x"0000" -- 4AC8
           ,x"4518" -- 4ACA
           ,x"6a00" -- 4ACC
           ,x"0000" -- 4ACE
           ,x"45f4" -- 4AD0
           ,x"2400" -- 4AD2
           ,x"0000" -- 4AD4
           ,x"4698" -- 4AD6
           ,x"9680" -- 4AD8
           ,x"0000" -- 4ADA
           ,x"475f" -- 4ADC
           ,x"5e10" -- 4ADE
           ,x"0000" -- 4AE0
           ,x"483b" -- 4AE2
           ,x"9aca" -- 4AE4
           ,x"0000" -- 4AE6
           ,x"ef88" -- 4AE8
           ,x"b4ec" -- 4AEA
           ,x"c22d" -- 4AEC
           ,x"0010" -- 4AEE
           ,x"9818" -- 4AF0
           ,x"80bc" -- 4AF2
           ,x"130c" -- 4AF4
           ,x"1a09" -- 4AF6
           ,x"9838" -- 4AF8
           ,x"c842" -- 4AFA
           ,x"1b06" -- 4AFC
           ,x"c088" -- 4AFE
           ,x"d038" -- 4B00
           ,x"16fe" -- 4B02
           ,x"04c0" -- 4B04
           ,x"d038" -- 4B06
           ,x"101f" -- 4B08
           ,x"8fbe" -- 4B0A
           ,x"0380" -- 4B0C
           ,x"05ce" -- 4B0E
           ,x"05ad" -- 4B10
           ,x"0010" -- 4B12
           ,x"04c5" -- 4B14
           ,x"06a0" -- 4B16
           ,x"b6d0" -- 4B18
           ,x"0282" -- 4B1A
           ,x"ee0c" -- 4B1C
           ,x"1a14" -- 4B1E
           ,x"0420" -- 4B20
           ,x"8d70" -- 4B22
           ,x"0016" -- 4B24
           ,x"ef88" -- 4B26
           ,x"b514" -- 4B28
           ,x"d818" -- 4B2A
           ,x"ede8" -- 4B2C
           ,x"1307" -- 4B2E
           ,x"9818" -- 4B30
           ,x"ab7f" -- 4B32
           ,x"1a03" -- 4B34
           ,x"9818" -- 4B36
           ,x"baa2" -- 4B38
           ,x"1a01" -- 4B3A
           ,x"05cb" -- 4B3C
           ,x"045b" -- 4B3E
           ,x"ef88" -- 4B40
           ,x"b544" -- 4B42
           ,x"06a0" -- 4B44
           ,x"b6ce" -- 4B46
           ,x"cb42" -- 4B48
           ,x"0004" -- 4B4A
           ,x"c800" -- 4B4C
           ,x"ede8" -- 4B4E
           ,x"c740" -- 4B50
           ,x"cb48" -- 4B52
           ,x"0010" -- 4B54
           ,x"0380" -- 4B56
           ,x"ef88" -- 4B58
           ,x"b55c" -- 4B5A
           ,x"c80b" -- 4B5C
           ,x"ed2c" -- 4B5E
           ,x"06a0" -- 4B60
           ,x"b6ce" -- 4B62
           ,x"06a0" -- 4B64
           ,x"bbd6" -- 4B66
           ,x"c320" -- 4B68
           ,x"ed2c" -- 4B6A
           ,x"c701" -- 4B6C
           ,x"10ee" -- 4B6E
           ,x"0420" -- 4B70
           ,x"8d70" -- 4B72
           ,x"0026" -- 4B74
           ,x"cd85" -- 4B76
           ,x"c106" -- 4B78
           ,x"c0e0" -- 4B7A
           ,x"ed0c" -- 4B7C
           ,x"0960" -- 4B7E
           ,x"a0c0" -- 4B80
           ,x"cdb3" -- 4B82
           ,x"13f5" -- 4B84
           ,x"c053" -- 4B86
           ,x"132d" -- 4B88
           ,x"c0e0" -- 4B8A
           ,x"edd6" -- 4B8C
           ,x"cdb3" -- 4B8E
           ,x"cdb3" -- 4B90
           ,x"cd93" -- 4B92
           ,x"0223" -- 4B94
           ,x"fffc" -- 4B96
           ,x"0705" -- 4B98
           ,x"9838" -- 4B9A
           ,x"ad1f" -- 4B9C
           ,x"1303" -- 4B9E
           ,x"0608" -- 4BA0
           ,x"04c5" -- 4BA2
           ,x"0701" -- 4BA4
           ,x"cd81" -- 4BA6
           ,x"cd83" -- 4BA8
           ,x"cd84" -- 4BAA
           ,x"06a0" -- 4BAC
           ,x"b6dc" -- 4BAE
           ,x"0646" -- 4BB0
           ,x"c116" -- 4BB2
           ,x"0646" -- 4BB4
           ,x"c0d6" -- 4BB6
           ,x"0646" -- 4BB8
           ,x"c056" -- 4BBA
           ,x"ccc6" -- 4BBC
           ,x"cdb2" -- 4BBE
           ,x"cdb2" -- 4BC0
           ,x"cd92" -- 4BC2
           ,x"0581" -- 4BC4
           ,x"1309" -- 4BC6
           ,x"0641" -- 4BC8
           ,x"1309" -- 4BCA
           ,x"0705" -- 4BCC
           ,x"0280" -- 4BCE
           ,x"3f00" -- 4BD0
           ,x"13e9" -- 4BD2
           ,x"0420" -- 4BD4
           ,x"8d70" -- 4BD6
           ,x"0025" -- 4BD8
           ,x"0608" -- 4BDA
           ,x"1003" -- 4BDC
           ,x"0280" -- 4BDE
           ,x"4b00" -- 4BE0
           ,x"16f8" -- 4BE2
           ,x"cd84" -- 4BE4
           ,x"cd88" -- 4BE6
           ,x"c214" -- 4BE8
           ,x"0705" -- 4BEA
           ,x"06a0" -- 4BEC
           ,x"b6dc" -- 4BEE
           ,x"0646" -- 4BF0
           ,x"c216" -- 4BF2
           ,x"0646" -- 4BF4
           ,x"c196" -- 4BF6
           ,x"c106" -- 4BF8
           ,x"05c4" -- 4BFA
           ,x"c0e0" -- 4BFC
           ,x"edd6" -- 4BFE
           ,x"ccf4" -- 4C00
           ,x"ccf4" -- 4C02
           ,x"c4d4" -- 4C04
           ,x"1052" -- 4C06
           ,x"9818" -- 4C08
           ,x"80bc" -- 4C0A
           ,x"130b" -- 4C0C
           ,x"1a09" -- 4C0E
           ,x"9818" -- 4C10
           ,x"c842" -- 4C12
           ,x"1b06" -- 4C14
           ,x"0588" -- 4C16
           ,x"c088" -- 4C18
           ,x"d038" -- 4C1A
           ,x"16fe" -- 4C1C
           ,x"d038" -- 4C1E
           ,x"05cb" -- 4C20
           ,x"045b" -- 4C22
           ,x"0588" -- 4C24
           ,x"05cb" -- 4C26
           ,x"04c5" -- 4C28
           ,x"0460" -- 4C2A
           ,x"b6dc" -- 4C2C
           ,x"cd85" -- 4C2E
           ,x"cd80" -- 4C30
           ,x"0201" -- 4C32
           ,x"0001" -- 4C34
           ,x"9838" -- 4C36
           ,x"ad1f" -- 4C38
           ,x"1306" -- 4C3A
           ,x"04c5" -- 4C3C
           ,x"0608" -- 4C3E
           ,x"06a0" -- 4C40
           ,x"b6dc" -- 4C42
           ,x"0608" -- 4C44
           ,x"1029" -- 4C46
           ,x"06a0" -- 4C48
           ,x"b608" -- 4C4A
           ,x"1009" -- 4C4C
           ,x"cd82" -- 4C4E
           ,x"0280" -- 4C50
           ,x"3f00" -- 4C52
           ,x"161d" -- 4C54
           ,x"06a0" -- 4C56
           ,x"b608" -- 4C58
           ,x"10bc" -- 4C5A
           ,x"c042" -- 4C5C
           ,x"1018" -- 4C5E
           ,x"0705" -- 4C60
           ,x"06a0" -- 4C62
           ,x"b6dc" -- 4C64
           ,x"0280" -- 4C66
           ,x"4b00" -- 4C68
           ,x"1317" -- 4C6A
           ,x"0280" -- 4C6C
           ,x"3f00" -- 4C6E
           ,x"16b1" -- 4C70
           ,x"8182" -- 4C72
           ,x"1a07" -- 4C74
           ,x"020b" -- 4C76
           ,x"edf2" -- 4C78
           ,x"c142" -- 4C7A
           ,x"c08b" -- 4C7C
           ,x"cef5" -- 4C7E
           ,x"cef5" -- 4C80
           ,x"c6d5" -- 4C82
           ,x"cd82" -- 4C84
           ,x"0705" -- 4C86
           ,x"06a0" -- 4C88
           ,x"b6dc" -- 4C8A
           ,x"06a0" -- 4C8C
           ,x"bbd6" -- 4C8E
           ,x"0646" -- 4C90
           ,x"c096" -- 4C92
           ,x"0280" -- 4C94
           ,x"4b00" -- 4C96
           ,x"169d" -- 4C98
           ,x"0646" -- 4C9A
           ,x"c0d6" -- 4C9C
           ,x"0973" -- 4C9E
           ,x"c2e3" -- 4CA0
           ,x"b8f6" -- 4CA2
           ,x"1309" -- 4CA4
           ,x"0420" -- 4CA6
           ,x"be74" -- 4CA8
           ,x"069b" -- 4CAA
           ,x"0646" -- 4CAC
           ,x"c156" -- 4CAE
           ,x"cdb2" -- 4CB0
           ,x"cdb2" -- 4CB2
           ,x"cd92" -- 4CB4
           ,x"106e" -- 4CB6
           ,x"0420" -- 4CB8
           ,x"8d70" -- 4CBA
           ,x"ffff" -- 4CBC
           ,x"0202" -- 4CBE
           ,x"ef68" -- 4CC0
           ,x"10f4" -- 4CC2
           ,x"0420" -- 4CC4
           ,x"c588" -- 4CC6
           ,x"0202" -- 4CC8
           ,x"ef68" -- 4CCA
           ,x"10f1" -- 4CCC
           ,x"0705" -- 4CCE
           ,x"c22d" -- 4CD0
           ,x"0010" -- 4CD2
           ,x"0206" -- 4CD4
           ,x"ee0c" -- 4CD6
           ,x"0207" -- 4CD8
           ,x"eea0" -- 4CDA
           ,x"cd8b" -- 4CDC
           ,x"04f6" -- 4CDE
           ,x"04c0" -- 4CE0
           ,x"d140" -- 4CE2
           ,x"0607" -- 4CE4
           ,x"d5c0" -- 4CE6
           ,x"81c6" -- 4CE8
           ,x"145b" -- 4CEA
           ,x"d038" -- 4CEC
           ,x"137e" -- 4CEE
           ,x"0280" -- 4CF0
           ,x"6f00" -- 4CF2
           ,x"1b24" -- 4CF4
           ,x"130f" -- 4CF6
           ,x"0280" -- 4CF8
           ,x"6200" -- 4CFA
           ,x"1413" -- 4CFC
           ,x"0280" -- 4CFE
           ,x"4c00" -- 4D00
           ,x"1b6c" -- 4D02
           ,x"13ef" -- 4D04
           ,x"0280" -- 4D06
           ,x"3800" -- 4D08
           ,x"1470" -- 4D0A
           ,x"0280" -- 4D0C
           ,x"1b00" -- 4D0E
           ,x"148e" -- 4D10
           ,x"0460" -- 4D12
           ,x"b576" -- 4D14
           ,x"ddb8" -- 4D16
           ,x"ddb8" -- 4D18
           ,x"ddb8" -- 4D1A
           ,x"ddb8" -- 4D1C
           ,x"ddb8" -- 4D1E
           ,x"ddb8" -- 4D20
           ,x"1038" -- 4D22
           ,x"0280" -- 4D24
           ,x"6d00" -- 4D26
           ,x"142e" -- 4D28
           ,x"06c0" -- 4D2A
           ,x"0220" -- 4D2C
           ,x"ff9d" -- 4D2E
           ,x"102e" -- 4D30
           ,x"0420" -- 4D32
           ,x"8d70" -- 4D34
           ,x"000a" -- 4D36
           ,x"0200" -- 4D38
           ,x"6100" -- 4D3A
           ,x"10d3" -- 4D3C
           ,x"0280" -- 4D3E
           ,x"7300" -- 4D40
           ,x"13c0" -- 4D42
           ,x"c060" -- 4D44
           ,x"edd4" -- 4D46
           ,x"0970" -- 4D48
           ,x"a040" -- 4D4A
           ,x"c061" -- 4D4C
           ,x"ff20" -- 4D4E
           ,x"1116" -- 4D50
           ,x"c060" -- 4D52
           ,x"edd6" -- 4D54
           ,x"a040" -- 4D56
           ,x"c021" -- 4D58
           ,x"ff20" -- 4D5A
           ,x"161c" -- 4D5C
           ,x"06c5" -- 4D5E
           ,x"d145" -- 4D60
           ,x"06c5" -- 4D62
           ,x"160d" -- 4D64
           ,x"c020" -- 4D66
           ,x"edda" -- 4D68
           ,x"0220" -- 4D6A
           ,x"fffa" -- 4D6C
           ,x"8800" -- 4D6E
           ,x"edd8" -- 4D70
           ,x"1adf" -- 4D72
           ,x"c840" -- 4D74
           ,x"ff20" -- 4D76
           ,x"c800" -- 4D78
           ,x"edda" -- 4D7A
           ,x"100c" -- 4D7C
           ,x"106e" -- 4D7E
           ,x"0420" -- 4D80
           ,x"8d70" -- 4D82
           ,x"0028" -- 4D84
           ,x"d038" -- 4D86
           ,x"06c0" -- 4D88
           ,x"d038" -- 4D8A
           ,x"06c0" -- 4D8C
           ,x"04f6" -- 4D8E
           ,x"cd80" -- 4D90
           ,x"04f6" -- 4D92
           ,x"0700" -- 4D94
           ,x"cd80" -- 4D96
           ,x"04c0" -- 4D98
           ,x"d160" -- 4D9A
           ,x"aa66" -- 4D9C
           ,x"81c6" -- 4D9E
           ,x"1aa5" -- 4DA0
           ,x"0420" -- 4DA2
           ,x"8d70" -- 4DA4
           ,x"001b" -- 4DA6
           ,x"0280" -- 4DA8
           ,x"5d00" -- 4DAA
           ,x"139f" -- 4DAC
           ,x"0280" -- 4DAE
           ,x"5c00" -- 4DB0
           ,x"13c2" -- 4DB2
           ,x"0280" -- 4DB4
           ,x"5200" -- 4DB6
           ,x"1395" -- 4DB8
           ,x"0280" -- 4DBA
           ,x"5300" -- 4DBC
           ,x"1392" -- 4DBE
           ,x"0420" -- 4DC0
           ,x"8d70" -- 4DC2
           ,x"0001" -- 4DC4
           ,x"0280" -- 4DC6
           ,x"4d00" -- 4DC8
           ,x"1612" -- 4DCA
           ,x"9817" -- 4DCC
           ,x"baa2" -- 4DCE
           ,x"160f" -- 4DD0
           ,x"0587" -- 4DD2
           ,x"108b" -- 4DD4
           ,x"d057" -- 4DD6
           ,x"16f9" -- 4DD8
           ,x"1008" -- 4DDA
           ,x"d045" -- 4DDC
           ,x"13e4" -- 4DDE
           ,x"0280" -- 4DE0
           ,x"4d00" -- 4DE2
           ,x"13f8" -- 4DE4
           ,x"0245" -- 4DE6
           ,x"00ff" -- 4DE8
           ,x"1602" -- 4DEA
           ,x"04c5" -- 4DEC
           ,x"04c0" -- 4DEE
           ,x"d057" -- 4DF0
           ,x"c100" -- 4DF2
           ,x"0244" -- 4DF4
           ,x"fe00" -- 4DF6
           ,x"9044" -- 4DF8
           ,x"1ba0" -- 4DFA
           ,x"d0f7" -- 4DFC
           ,x"131c" -- 4DFE
           ,x"0973" -- 4E00
           ,x"c2e3" -- 4E02
           ,x"b85a" -- 4E04
           ,x"0646" -- 4E06
           ,x"c056" -- 4E08
           ,x"13da" -- 4E0A
           ,x"0596" -- 4E0C
           ,x"1603" -- 4E0E
           ,x"0226" -- 4E10
           ,x"fffa" -- 4E12
           ,x"c046" -- 4E14
           ,x"22e0" -- 4E16
           ,x"b920" -- 4E18
           ,x"1308" -- 4E1A
           ,x"0646" -- 4E1C
           ,x"c096" -- 4E1E
           ,x"13cf" -- 4E20
           ,x"0596" -- 4E22
           ,x"1603" -- 4E24
           ,x"0226" -- 4E26
           ,x"fffa" -- 4E28
           ,x"c086" -- 4E2A
           ,x"069b" -- 4E2C
           ,x"cdb2" -- 4E2E
           ,x"cdb2" -- 4E30
           ,x"cd92" -- 4E32
           ,x"0736" -- 4E34
           ,x"10c7" -- 4E36
           ,x"d028" -- 4E38
           ,x"ffff" -- 4E3A
           ,x"0646" -- 4E3C
           ,x"c096" -- 4E3E
           ,x"13bf" -- 4E40
           ,x"0596" -- 4E42
           ,x"1603" -- 4E44
           ,x"0226" -- 4E46
           ,x"fffa" -- 4E48
           ,x"c086" -- 4E4A
           ,x"0226" -- 4E4C
           ,x"fffc" -- 4E4E
           ,x"c2d6" -- 4E50
           ,x"c066" -- 4E52
           ,x"0002" -- 4E54
           ,x"16b4" -- 4E56
           ,x"045b" -- 4E58
           ,x"109f" -- 4E5A
           ,x"c060" -- 4E5C
           ,x"edd6" -- 4E5E
           ,x"a040" -- 4E60
           ,x"c121" -- 4E62
           ,x"ff20" -- 4E64
           ,x"1341" -- 4E66
           ,x"cd85" -- 4E68
           ,x"04f6" -- 4E6A
           ,x"cd84" -- 4E6C
           ,x"0705" -- 4E6E
           ,x"06a0" -- 4E70
           ,x"b6dc" -- 4E72
           ,x"06a0" -- 4E74
           ,x"bbd6" -- 4E76
           ,x"0646" -- 4E78
           ,x"c116" -- 4E7A
           ,x"0646" -- 4E7C
           ,x"8d01" -- 4E7E
           ,x"1b2e" -- 4E80
           ,x"c174" -- 4E82
           ,x"0285" -- 4E84
           ,x"ffff" -- 4E86
           ,x"1308" -- 4E88
           ,x"3845" -- 4E8A
           ,x"ad82" -- 4E8C
           ,x"0280" -- 4E8E
           ,x"3f00" -- 4E90
           ,x"13ec" -- 4E92
           ,x"0420" -- 4E94
           ,x"8d70" -- 4E96
           ,x"0012" -- 4E98
           ,x"a056" -- 4E9A
           ,x"3860" -- 4E9C
           ,x"b92a" -- 4E9E
           ,x"a084" -- 4EA0
           ,x"0646" -- 4EA2
           ,x"c156" -- 4EA4
           ,x"cd82" -- 4EA6
           ,x"0280" -- 4EA8
           ,x"4b00" -- 4EAA
           ,x"13d6" -- 4EAC
           ,x"0280" -- 4EAE
           ,x"4000" -- 4EB0
           ,x"1618" -- 4EB2
           ,x"cd85" -- 4EB4
           ,x"0705" -- 4EB6
           ,x"06a0" -- 4EB8
           ,x"b6dc" -- 4EBA
           ,x"06a0" -- 4EBC
           ,x"bbd6" -- 4EBE
           ,x"0280" -- 4EC0
           ,x"4b00" -- 4EC2
           ,x"1615" -- 4EC4
           ,x"0646" -- 4EC6
           ,x"c156" -- 4EC8
           ,x"0646" -- 4ECA
           ,x"c016" -- 4ECC
           ,x"0601" -- 4ECE
           ,x"1106" -- 4ED0
           ,x"a001" -- 4ED2
           ,x"8800" -- 4ED4
           ,x"ed04" -- 4ED6
           ,x"1402" -- 4ED8
           ,x"0460" -- 4EDA
           ,x"b796" -- 4EDC
           ,x"0420" -- 4EDE
           ,x"8d70" -- 4EE0
           ,x"0011" -- 4EE2
           ,x"0420" -- 4EE4
           ,x"8d70" -- 4EE6
           ,x"0013" -- 4EE8
           ,x"0420" -- 4EEA
           ,x"8d70" -- 4EEC
           ,x"0027" -- 4EEE
           ,x"0420" -- 4EF0
           ,x"8d70" -- 4EF2
           ,x"0025" -- 4EF4
           ,x"a330" -- 4EF6
           ,x"994e" -- 4EF8
           ,x"a312" -- 4EFA
           ,x"9960" -- 4EFC
           ,x"a347" -- 4EFE
           ,x"9973" -- 4F00
           ,x"9956" -- 4F02
           ,x"ba46" -- 4F04
           ,x"ba46" -- 4F06
           ,x"ba46" -- 4F08
           ,x"ba46" -- 4F0A
           ,x"ba46" -- 4F0C
           ,x"ba46" -- 4F0E
           ,x"ba46" -- 4F10
           ,x"b9be" -- 4F12
           ,x"b98e" -- 4F14
           ,x"ba04" -- 4F16
           ,x"b9ce" -- 4F18
           ,x"c53a" -- 4F1A
           ,x"ba85" -- 4F1C
           ,x"0000" -- 4F1E
           ,x"0001" -- 4F20
           ,x"0004" -- 4F22
           ,x"0005" -- 4F24
           ,x"0002" -- 4F26
           ,x"0003" -- 4F28
           ,x"0006" -- 4F2A
           ,x"9440" -- 4F2C
           ,x"9a4c" -- 4F2E
           ,x"99b6" -- 4F30
           ,x"8778" -- 4F32
           ,x"c5a0" -- 4F34
           ,x"baaa" -- 4F36
           ,x"9486" -- 4F38
           ,x"940a" -- 4F3A
           ,x"c1e0" -- 4F3C
           ,x"946c" -- 4F3E
           ,x"c5ba" -- 4F40
           ,x"c67c" -- 4F42
           ,x"93e4" -- 4F44
           ,x"a246" -- 4F46
           ,x"a168" -- 4F48
           ,x"bfde" -- 4F4A
           ,x"8fa6" -- 4F4C
           ,x"8f7c" -- 4F4E
           ,x"99a2" -- 4F50
           ,x"9a3a" -- 4F52
           ,x"8f2e" -- 4F54
           ,x"8f20" -- 4F56
           ,x"8efc" -- 4F58
           ,x"8a84" -- 4F5A
           ,x"94d0" -- 4F5C
           ,x"0000" -- 4F5E
           ,x"0000" -- 4F60
           ,x"0000" -- 4F62
           ,x"0000" -- 4F64
           ,x"c811" -- 4F66
           ,x"ef60" -- 4F68
           ,x"c821" -- 4F6A
           ,x"0002" -- 4F6C
           ,x"ef62" -- 4F6E
           ,x"c821" -- 4F70
           ,x"0004" -- 4F72
           ,x"ef64" -- 4F74
           ,x"c802" -- 4F76
           ,x"ef7e" -- 4F78
           ,x"0420" -- 4F7A
           ,x"bc3e" -- 4F7C
           ,x"c0f1" -- 4F7E
           ,x"160d" -- 4F80
           ,x"c0f2" -- 4F82
           ,x"160b" -- 4F84
           ,x"c0d1" -- 4F86
           ,x"c052" -- 4F88
           ,x"046b" -- 4F8A
           ,x"0004" -- 4F8C
           ,x"c28b" -- 4F8E
           ,x"06a0" -- 4F90
           ,x"b966" -- 4F92
           ,x"ef68" -- 4F94
           ,x"bc5c" -- 4F96
           ,x"a043" -- 4F98
           ,x"190a" -- 4F9A
           ,x"0420" -- 4F9C
           ,x"b9ba" -- 4F9E
           ,x"0420" -- 4FA0
           ,x"bd1a" -- 4FA2
           ,x"c820" -- 4FA4
           ,x"8012" -- 4FA6
           ,x"ef7e" -- 4FA8
           ,x"041b" -- 4FAA
           ,x"1003" -- 4FAC
           ,x"0501" -- 4FAE
           ,x"c801" -- 4FB0
           ,x"ef6a" -- 4FB2
           ,x"0202" -- 4FB4
           ,x"ef68" -- 4FB6
           ,x"045a" -- 4FB8
           ,x"ef60" -- 4FBA
           ,x"bd1e" -- 4FBC
           ,x"c28b" -- 4FBE
           ,x"06a0" -- 4FC0
           ,x"b966" -- 4FC2
           ,x"ef68" -- 4FC4
           ,x"bc52" -- 4FC6
           ,x"6043" -- 4FC8
           ,x"19f2" -- 4FCA
           ,x"10e7" -- 4FCC
           ,x"c28b" -- 4FCE
           ,x"06a0" -- 4FD0
           ,x"b966" -- 4FD2
           ,x"ef68" -- 4FD4
           ,x"bd88" -- 4FD6
           ,x"c0c3" -- 4FD8
           ,x"1108" -- 4FDA
           ,x"c041" -- 4FDC
           ,x"110b" -- 4FDE
           ,x"3843" -- 4FE0
           ,x"c041" -- 4FE2
           ,x"16db" -- 4FE4
           ,x"c042" -- 4FE6
           ,x"11d9" -- 4FE8
           ,x"10e2" -- 4FEA
           ,x"0503" -- 4FEC
           ,x"c041" -- 4FEE
           ,x"1503" -- 4FF0
           ,x"0501" -- 4FF2
           ,x"10f5" -- 4FF4
           ,x"0501" -- 4FF6
           ,x"3843" -- 4FF8
           ,x"c041" -- 4FFA
           ,x"16cf" -- 4FFC
           ,x"c042" -- 4FFE
           ,x"11cd" -- 5000
           ,x"10d5" -- 5002
           ,x"c28b" -- 5004
           ,x"06a0" -- 5006
           ,x"b966" -- 5008
           ,x"ef68" -- 500A
           ,x"beb0" -- 500C
           ,x"c0c3" -- 500E
           ,x"110a" -- 5010
           ,x"1316" -- 5012
           ,x"c081" -- 5014
           ,x"110c" -- 5016
           ,x"04c1" -- 5018
           ,x"3c43" -- 501A
           ,x"c082" -- 501C
           ,x"16be" -- 501E
           ,x"c041" -- 5020
           ,x"11bc" -- 5022
           ,x"10c5" -- 5024
           ,x"0503" -- 5026
           ,x"c081" -- 5028
           ,x"1503" -- 502A
           ,x"0502" -- 502C
           ,x"10f4" -- 502E
           ,x"0502" -- 5030
           ,x"04c1" -- 5032
           ,x"3c43" -- 5034
           ,x"c082" -- 5036
           ,x"16b1" -- 5038
           ,x"c041" -- 503A
           ,x"11af" -- 503C
           ,x"10b7" -- 503E
           ,x"0420" -- 5040
           ,x"8d70" -- 5042
           ,x"001c" -- 5044
           ,x"c123" -- 5046
           ,x"b874" -- 5048
           ,x"06a0" -- 504A
           ,x"b9be" -- 504C
           ,x"0203" -- 504E
           ,x"0004" -- 5050
           ,x"c104" -- 5052
           ,x"1609" -- 5054
           ,x"0584" -- 5056
           ,x"c052" -- 5058
           ,x"1306" -- 505A
           ,x"0241" -- 505C
           ,x"7f00" -- 505E
           ,x"0281" -- 5060
           ,x"3b00" -- 5062
           ,x"1a06" -- 5064
           ,x"1007" -- 5066
           ,x"c072" -- 5068
           ,x"1601" -- 506A
           ,x"c052" -- 506C
           ,x"1503" -- 506E
           ,x"1601" -- 5070
           ,x"0603" -- 5072
           ,x"0643" -- 5074
           ,x"0420" -- 5076
           ,x"be74" -- 5078
           ,x"2103" -- 507A
           ,x"160e" -- 507C
           ,x"05a0" -- 507E
           ,x"ef6a" -- 5080
           ,x"100b" -- 5082
           ,x"c801" -- 5084
           ,x"ef7e" -- 5086
           ,x"0420" -- 5088
           ,x"bc3e" -- 508A
           ,x"c051" -- 508C
           ,x"1303" -- 508E
           ,x"0420" -- 5090
           ,x"bd0c" -- 5092
           ,x"1002" -- 5094
           ,x"0520" -- 5096
           ,x"ef6a" -- 5098
           ,x"0202" -- 509A
           ,x"ef68" -- 509C
           ,x"0460" -- 509E
           ,x"b82e" -- 50A0
           ,x"4c00" -- 50A2
           ,x"0420" -- 50A4
           ,x"8d70" -- 50A6
           ,x"0021" -- 50A8
           ,x"c28b" -- 50AA
           ,x"06a0" -- 50AC
           ,x"c4d0" -- 50AE
           ,x"1366" -- 50B0
           ,x"c820" -- 50B2
           ,x"bb8e" -- 50B4
           ,x"ef7e" -- 50B6
           ,x"0420" -- 50B8
           ,x"bd84" -- 50BA
           ,x"06a0" -- 50BC
           ,x"c48c" -- 50BE
           ,x"0281" -- 50C0
           ,x"007d" -- 50C2
           ,x"15ef" -- 50C4
           ,x"c081" -- 50C6
           ,x"c820" -- 50C8
           ,x"bb90" -- 50CA
           ,x"ef7e" -- 50CC
           ,x"0420" -- 50CE
           ,x"bc4e" -- 50D0
           ,x"c820" -- 50D2
           ,x"8000" -- 50D4
           ,x"ef7e" -- 50D6
           ,x"0420" -- 50D8
           ,x"bc32" -- 50DA
           ,x"06a0" -- 50DC
           ,x"c4f4" -- 50DE
           ,x"bba2" -- 50E0
           ,x"c820" -- 50E2
           ,x"8000" -- 50E4
           ,x"ef7e" -- 50E6
           ,x"0420" -- 50E8
           ,x"bd84" -- 50EA
           ,x"c820" -- 50EC
           ,x"8000" -- 50EE
           ,x"ef7e" -- 50F0
           ,x"0420" -- 50F2
           ,x"bc32" -- 50F4
           ,x"06a0" -- 50F6
           ,x"c512" -- 50F8
           ,x"bbb6" -- 50FA
           ,x"c820" -- 50FC
           ,x"8012" -- 50FE
           ,x"ef7e" -- 5100
           ,x"0420" -- 5102
           ,x"bc32" -- 5104
           ,x"c820" -- 5106
           ,x"8000" -- 5108
           ,x"ef7e" -- 510A
           ,x"0420" -- 510C
           ,x"bc4e" -- 510E
           ,x"c820" -- 5110
           ,x"8002" -- 5112
           ,x"ef7e" -- 5114
           ,x"0420" -- 5116
           ,x"bc32" -- 5118
           ,x"c820" -- 511A
           ,x"8012" -- 511C
           ,x"ef7e" -- 511E
           ,x"0420" -- 5120
           ,x"bc3e" -- 5122
           ,x"c820" -- 5124
           ,x"8000" -- 5126
           ,x"ef7e" -- 5128
           ,x"0420" -- 512A
           ,x"bc4a" -- 512C
           ,x"c820" -- 512E
           ,x"8002" -- 5130
           ,x"ef7e" -- 5132
           ,x"0420" -- 5134
           ,x"beac" -- 5136
           ,x"c820" -- 5138
           ,x"bb94" -- 513A
           ,x"ef7e" -- 513C
           ,x"0420" -- 513E
           ,x"bd84" -- 5140
           ,x"c042" -- 5142
           ,x"0921" -- 5144
           ,x"06c1" -- 5146
           ,x"a801" -- 5148
           ,x"ef68" -- 514A
           ,x"c043" -- 514C
           ,x"0242" -- 514E
           ,x"0003" -- 5150
           ,x"1303" -- 5152
           ,x"c0c2" -- 5154
           ,x"06a0" -- 5156
           ,x"c18a" -- 5158
           ,x"c041" -- 515A
           ,x"1315" -- 515C
           ,x"c820" -- 515E
           ,x"8012" -- 5160
           ,x"ef7e" -- 5162
           ,x"0420" -- 5164
           ,x"bc32" -- 5166
           ,x"c820" -- 5168
           ,x"bb92" -- 516A
           ,x"ef7e" -- 516C
           ,x"0420" -- 516E
           ,x"bc3e" -- 5170
           ,x"c820" -- 5172
           ,x"8012" -- 5174
           ,x"ef7e" -- 5176
           ,x"0420" -- 5178
           ,x"beac" -- 517A
           ,x"1005" -- 517C
           ,x"c820" -- 517E
           ,x"bb92" -- 5180
           ,x"ef7e" -- 5182
           ,x"0420" -- 5184
           ,x"bc3e" -- 5186
           ,x"0202" -- 5188
           ,x"ef68" -- 518A
           ,x"045a" -- 518C
           ,x"bb96" -- 518E
           ,x"bb9c" -- 5190
           ,x"bbb8" -- 5192
           ,x"bbd0" -- 5194
           ,x"4117" -- 5196
           ,x"1547" -- 5198
           ,x"652c" -- 519A
           ,x"4080" -- 519C
           ,x"0000" -- 519E
           ,x"0000" -- 51A0
           ,x"0002" -- 51A2
           ,x"423c" -- 51A4
           ,x"9d67" -- 51A6
           ,x"06a2" -- 51A8
           ,x"4476" -- 51AA
           ,x"4ef8" -- 51AC
           ,x"c12a" -- 51AE
           ,x"461f" -- 51B0
           ,x"be80" -- 51B2
           ,x"58c1" -- 51B4
           ,x"0003" -- 51B6
           ,x"4110" -- 51B8
           ,x"0000" -- 51BA
           ,x"0000" -- 51BC
           ,x"436d" -- 51BE
           ,x"549a" -- 51C0
           ,x"5fe1" -- 51C2
           ,x"4550" -- 51C4
           ,x"02d2" -- 51C6
           ,x"6dcf" -- 51C8
           ,x"465b" -- 51CA
           ,x"9820" -- 51CC
           ,x"5c39" -- 51CE
           ,x"4116" -- 51D0
           ,x"a09e" -- 51D2
           ,x"667f" -- 51D4
           ,x"c072" -- 51D6
           ,x"1602" -- 51D8
           ,x"c052" -- 51DA
           ,x"045b" -- 51DC
           ,x"c802" -- 51DE
           ,x"ef7e" -- 51E0
           ,x"0660" -- 51E2
           ,x"ef7e" -- 51E4
           ,x"0420" -- 51E6
           ,x"bc3e" -- 51E8
           ,x"c081" -- 51EA
           ,x"0241" -- 51EC
           ,x"7f80" -- 51EE
           ,x"0281" -- 51F0
           ,x"4400" -- 51F2
           ,x"150d" -- 51F4
           ,x"c820" -- 51F6
           ,x"c83e" -- 51F8
           ,x"ef7e" -- 51FA
           ,x"0420" -- 51FC
           ,x"bf7c" -- 51FE
           ,x"c060" -- 5200
           ,x"ef6a" -- 5202
           ,x"0420" -- 5204
           ,x"be74" -- 5206
           ,x"0a12" -- 5208
           ,x"1701" -- 520A
           ,x"0501" -- 520C
           ,x"045b" -- 520E
           ,x"0420" -- 5210
           ,x"8d70" -- 5212
           ,x"001e" -- 5214
           ,x"c802" -- 5216
           ,x"ef7e" -- 5218
           ,x"0420" -- 521A
           ,x"bc3e" -- 521C
           ,x"c052" -- 521E
           ,x"1305" -- 5220
           ,x"c820" -- 5222
           ,x"c83e" -- 5224
           ,x"ef7e" -- 5226
           ,x"0420" -- 5228
           ,x"bf7c" -- 522A
           ,x"c060" -- 522C
           ,x"ef6a" -- 522E
           ,x"045b" -- 5230
           ,x"ef68" -- 5232
           ,x"bc36" -- 5234
           ,x"cec0" -- 5236
           ,x"cec1" -- 5238
           ,x"c6c2" -- 523A
           ,x"0380" -- 523C
           ,x"ef68" -- 523E
           ,x"bc42" -- 5240
           ,x"c03b" -- 5242
           ,x"c07b" -- 5244
           ,x"c09b" -- 5246
           ,x"0380" -- 5248
           ,x"ef68" -- 524A
           ,x"bc5c" -- 524C
           ,x"ef68" -- 524E
           ,x"bc52" -- 5250
           ,x"c13b" -- 5252
           ,x"13f9" -- 5254
           ,x"0224" -- 5256
           ,x"8000" -- 5258
           ,x"1002" -- 525A
           ,x"c13b" -- 525C
           ,x"13f4" -- 525E
           ,x"c000" -- 5260
           ,x"1602" -- 5262
           ,x"c004" -- 5264
           ,x"10ee" -- 5266
           ,x"c17b" -- 5268
           ,x"c19b" -- 526A
           ,x"d0c0" -- 526C
           ,x"d1c4" -- 526E
           ,x"7000" -- 5270
           ,x"7104" -- 5272
           ,x"0a13" -- 5274
           ,x"1702" -- 5276
           ,x"06a0" -- 5278
           ,x"bcfa" -- 527A
           ,x"0993" -- 527C
           ,x"0a17" -- 527E
           ,x"1708" -- 5280
           ,x"0506" -- 5282
           ,x"1604" -- 5284
           ,x"0505" -- 5286
           ,x"1603" -- 5288
           ,x"0504" -- 528A
           ,x"1002" -- 528C
           ,x"0545" -- 528E
           ,x"0544" -- 5290
           ,x"020a" -- 5292
           ,x"000a" -- 5294
           ,x"0997" -- 5296
           ,x"81c3" -- 5298
           ,x"131d" -- 529A
           ,x"1509" -- 529C
           ,x"06a0" -- 529E
           ,x"bf34" -- 52A0
           ,x"060a" -- 52A2
           ,x"16f9" -- 52A4
           ,x"c004" -- 52A6
           ,x"c045" -- 52A8
           ,x"c086" -- 52AA
           ,x"c0c7" -- 52AC
           ,x"100c" -- 52AE
           ,x"0946" -- 52B0
           ,x"c245" -- 52B2
           ,x"0ac9" -- 52B4
           ,x"a189" -- 52B6
           ,x"0945" -- 52B8
           ,x"c244" -- 52BA
           ,x"0ac9" -- 52BC
           ,x"a149" -- 52BE
           ,x"0844" -- 52C0
           ,x"0587" -- 52C2
           ,x"060a" -- 52C4
           ,x"16e8" -- 52C6
           ,x"c000" -- 52C8
           ,x"1559" -- 52CA
           ,x"06a0" -- 52CC
           ,x"bcfa" -- 52CE
           ,x"0223" -- 52D0
           ,x"0080" -- 52D2
           ,x"1054" -- 52D4
           ,x"06a0" -- 52D6
           ,x"bf54" -- 52D8
           ,x"1106" -- 52DA
           ,x"1509" -- 52DC
           ,x"c041" -- 52DE
           ,x"1607" -- 52E0
           ,x"c082" -- 52E2
           ,x"1605" -- 52E4
           ,x"104d" -- 52E6
           ,x"06a0" -- 52E8
           ,x"bcfa" -- 52EA
           ,x"0263" -- 52EC
           ,x"0080" -- 52EE
           ,x"d000" -- 52F0
           ,x"1334" -- 52F2
           ,x"06a0" -- 52F4
           ,x"bf34" -- 52F6
           ,x"1031" -- 52F8
           ,x"0502" -- 52FA
           ,x"1604" -- 52FC
           ,x"0501" -- 52FE
           ,x"1603" -- 5300
           ,x"0500" -- 5302
           ,x"045b" -- 5304
           ,x"0541" -- 5306
           ,x"0540" -- 5308
           ,x"045b" -- 530A
           ,x"ef68" -- 530C
           ,x"bd10" -- 530E
           ,x"c000" -- 5310
           ,x"1302" -- 5312
           ,x"0220" -- 5314
           ,x"8000" -- 5316
           ,x"0380" -- 5318
           ,x"ef68" -- 531A
           ,x"bd1e" -- 531C
           ,x"c000" -- 531E
           ,x"1630" -- 5320
           ,x"0203" -- 5322
           ,x"0044" -- 5324
           ,x"04c2" -- 5326
           ,x"c041" -- 5328
           ,x"1504" -- 532A
           ,x"1330" -- 532C
           ,x"0501" -- 532E
           ,x"0203" -- 5330
           ,x"00c4" -- 5332
           ,x"d001" -- 5334
           ,x"1303" -- 5336
           ,x"06c0" -- 5338
           ,x"0a81" -- 533A
           ,x"100f" -- 533C
           ,x"c001" -- 533E
           ,x"04c1" -- 5340
           ,x"0643" -- 5342
           ,x"100b" -- 5344
           ,x"ef68" -- 5346
           ,x"bd4a" -- 5348
           ,x"04c3" -- 534A
           ,x"d0c0" -- 534C
           ,x"6003" -- 534E
           ,x"1604" -- 5350
           ,x"c041" -- 5352
           ,x"1602" -- 5354
           ,x"c082" -- 5356
           ,x"1314" -- 5358
           ,x"06c3" -- 535A
           ,x"2420" -- 535C
           ,x"c848" -- 535E
           ,x"160e" -- 5360
           ,x"24e0" -- 5362
           ,x"c84a" -- 5364
           ,x"1313" -- 5366
           ,x"0603" -- 5368
           ,x"0a40" -- 536A
           ,x"c241" -- 536C
           ,x"09c9" -- 536E
           ,x"a009" -- 5370
           ,x"0a41" -- 5372
           ,x"c242" -- 5374
           ,x"09c9" -- 5376
           ,x"a049" -- 5378
           ,x"0a42" -- 537A
           ,x"10ef" -- 537C
           ,x"06c3" -- 537E
           ,x"d003" -- 5380
           ,x"0380" -- 5382
           ,x"ef68" -- 5384
           ,x"bd88" -- 5386
           ,x"c000" -- 5388
           ,x"1376" -- 538A
           ,x"c13b" -- 538C
           ,x"1374" -- 538E
           ,x"c17b" -- 5390
           ,x"c19b" -- 5392
           ,x"06a0" -- 5394
           ,x"be80" -- 5396
           ,x"a0c7" -- 5398
           ,x"ffc0" -- 539A
           ,x"c286" -- 539C
           ,x"3a82" -- 539E
           ,x"c206" -- 53A0
           ,x"3a01" -- 53A2
           ,x"3980" -- 53A4
           ,x"a289" -- 53A6
           ,x"1701" -- 53A8
           ,x"0588" -- 53AA
           ,x"a207" -- 53AC
           ,x"1701" -- 53AE
           ,x"0586" -- 53B0
           ,x"c248" -- 53B2
           ,x"c206" -- 53B4
           ,x"c185" -- 53B6
           ,x"3982" -- 53B8
           ,x"a287" -- 53BA
           ,x"1701" -- 53BC
           ,x"0586" -- 53BE
           ,x"a246" -- 53C0
           ,x"1701" -- 53C2
           ,x"0588" -- 53C4
           ,x"c289" -- 53C6
           ,x"c248" -- 53C8
           ,x"c1c5" -- 53CA
           ,x"39c1" -- 53CC
           ,x"3940" -- 53CE
           ,x"a288" -- 53D0
           ,x"04c8" -- 53D2
           ,x"1701" -- 53D4
           ,x"0587" -- 53D6
           ,x"a247" -- 53D8
           ,x"1701" -- 53DA
           ,x"0588" -- 53DC
           ,x"a246" -- 53DE
           ,x"1701" -- 53E0
           ,x"0588" -- 53E2
           ,x"04c7" -- 53E4
           ,x"a205" -- 53E6
           ,x"1701" -- 53E8
           ,x"0587" -- 53EA
           ,x"c144" -- 53EC
           ,x"3942" -- 53EE
           ,x"a286" -- 53F0
           ,x"1705" -- 53F2
           ,x"0589" -- 53F4
           ,x"1703" -- 53F6
           ,x"0588" -- 53F8
           ,x"1701" -- 53FA
           ,x"0587" -- 53FC
           ,x"a245" -- 53FE
           ,x"1703" -- 5400
           ,x"0588" -- 5402
           ,x"1701" -- 5404
           ,x"0587" -- 5406
           ,x"c144" -- 5408
           ,x"3941" -- 540A
           ,x"a246" -- 540C
           ,x"1703" -- 540E
           ,x"0588" -- 5410
           ,x"1701" -- 5412
           ,x"0587" -- 5414
           ,x"a205" -- 5416
           ,x"1701" -- 5418
           ,x"0587" -- 541A
           ,x"3900" -- 541C
           ,x"a205" -- 541E
           ,x"1701" -- 5420
           ,x"0587" -- 5422
           ,x"a1c4" -- 5424
           ,x"d1c8" -- 5426
           ,x"06c7" -- 5428
           ,x"d209" -- 542A
           ,x"06c8" -- 542C
           ,x"d24a" -- 542E
           ,x"06c9" -- 5430
           ,x"06ca" -- 5432
           ,x"c007" -- 5434
           ,x"c048" -- 5436
           ,x"c089" -- 5438
           ,x"2420" -- 543A
           ,x"c848" -- 543C
           ,x"1611" -- 543E
           ,x"24e0" -- 5440
           ,x"c84a" -- 5442
           ,x"1319" -- 5444
           ,x"0603" -- 5446
           ,x"0a40" -- 5448
           ,x"c241" -- 544A
           ,x"09c9" -- 544C
           ,x"a009" -- 544E
           ,x"0a41" -- 5450
           ,x"c242" -- 5452
           ,x"09c9" -- 5454
           ,x"a049" -- 5456
           ,x"0a42" -- 5458
           ,x"c24a" -- 545A
           ,x"09c9" -- 545C
           ,x"a089" -- 545E
           ,x"0a4a" -- 5460
           ,x"0a1a" -- 5462
           ,x"178c" -- 5464
           ,x"0582" -- 5466
           ,x"178a" -- 5468
           ,x"0581" -- 546A
           ,x"1788" -- 546C
           ,x"0580" -- 546E
           ,x"0460" -- 5470
           ,x"bcf0" -- 5472
           ,x"ef68" -- 5474
           ,x"be78" -- 5476
           ,x"04c0" -- 5478
           ,x"04c1" -- 547A
           ,x"04c2" -- 547C
           ,x"0380" -- 547E
           ,x"d0c0" -- 5480
           ,x"d1c4" -- 5482
           ,x"7000" -- 5484
           ,x"7104" -- 5486
           ,x"c207" -- 5488
           ,x"2a03" -- 548A
           ,x"06c3" -- 548C
           ,x"0243" -- 548E
           ,x"007f" -- 5490
           ,x"06c7" -- 5492
           ,x"0247" -- 5494
           ,x"007f" -- 5496
           ,x"04bb" -- 5498
           ,x"a0fb" -- 549A
           ,x"24e0" -- 549C
           ,x"aa66" -- 549E
           ,x"1646" -- 54A0
           ,x"0a18" -- 54A2
           ,x"1702" -- 54A4
           ,x"0223" -- 54A6
           ,x"0080" -- 54A8
           ,x"045b" -- 54AA
           ,x"ef68" -- 54AC
           ,x"beb0" -- 54AE
           ,x"c000" -- 54B0
           ,x"13e2" -- 54B2
           ,x"c13b" -- 54B4
           ,x"1338" -- 54B6
           ,x"c17b" -- 54B8
           ,x"c19b" -- 54BA
           ,x"06a0" -- 54BC
           ,x"be80" -- 54BE
           ,x"60c7" -- 54C0
           ,x"0040" -- 54C2
           ,x"8100" -- 54C4
           ,x"110a" -- 54C6
           ,x"0583" -- 54C8
           ,x"0a44" -- 54CA
           ,x"c245" -- 54CC
           ,x"09c9" -- 54CE
           ,x"a109" -- 54D0
           ,x"0a45" -- 54D2
           ,x"c246" -- 54D4
           ,x"09c9" -- 54D6
           ,x"a149" -- 54D8
           ,x"0a46" -- 54DA
           ,x"04c7" -- 54DC
           ,x"04c8" -- 54DE
           ,x"04c9" -- 54E0
           ,x"020a" -- 54E2
           ,x"0028" -- 54E4
           ,x"0a10" -- 54E6
           ,x"0a11" -- 54E8
           ,x"1701" -- 54EA
           ,x"0580" -- 54EC
           ,x"0a12" -- 54EE
           ,x"1701" -- 54F0
           ,x"0581" -- 54F2
           ,x"0a17" -- 54F4
           ,x"0a18" -- 54F6
           ,x"1701" -- 54F8
           ,x"0587" -- 54FA
           ,x"0a19" -- 54FC
           ,x"1701" -- 54FE
           ,x"0588" -- 5500
           ,x"8100" -- 5502
           ,x"1a09" -- 5504
           ,x"1b05" -- 5506
           ,x"8141" -- 5508
           ,x"1a06" -- 550A
           ,x"1b02" -- 550C
           ,x"8182" -- 550E
           ,x"1a03" -- 5510
           ,x"06a0" -- 5512
           ,x"bf68" -- 5514
           ,x"0589" -- 5516
           ,x"060a" -- 5518
           ,x"16e5" -- 551A
           ,x"0a10" -- 551C
           ,x"8100" -- 551E
           ,x"1a89" -- 5520
           ,x"020a" -- 5522
           ,x"8000" -- 5524
           ,x"1086" -- 5526
           ,x"0420" -- 5528
           ,x"8d70" -- 552A
           ,x"001c" -- 552C
           ,x"0420" -- 552E
           ,x"8d70" -- 5530
           ,x"001d" -- 5532
           ,x"0942" -- 5534
           ,x"c241" -- 5536
           ,x"0ac9" -- 5538
           ,x"a089" -- 553A
           ,x"0941" -- 553C
           ,x"c240" -- 553E
           ,x"0ac9" -- 5540
           ,x"a049" -- 5542
           ,x"0840" -- 5544
           ,x"c243" -- 5546
           ,x"0583" -- 5548
           ,x"2a43" -- 554A
           ,x"0249" -- 554C
           ,x"0080" -- 554E
           ,x"16ee" -- 5550
           ,x"045b" -- 5552
           ,x"a086" -- 5554
           ,x"1703" -- 5556
           ,x"0581" -- 5558
           ,x"1701" -- 555A
           ,x"0580" -- 555C
           ,x"a045" -- 555E
           ,x"1701" -- 5560
           ,x"0580" -- 5562
           ,x"a004" -- 5564
           ,x"045b" -- 5566
           ,x"6086" -- 5568
           ,x"1803" -- 556A
           ,x"0601" -- 556C
           ,x"1801" -- 556E
           ,x"0600" -- 5570
           ,x"6045" -- 5572
           ,x"1801" -- 5574
           ,x"0600" -- 5576
           ,x"6004" -- 5578
           ,x"045b" -- 557A
           ,x"ef68" -- 557C
           ,x"bf80" -- 557E
           ,x"c11b" -- 5580
           ,x"04c3" -- 5582
           ,x"c200" -- 5584
           ,x"d1c8" -- 5586
           ,x"0247" -- 5588
           ,x"7f00" -- 558A
           ,x"61c4" -- 558C
           ,x"130b" -- 558E
           ,x"d003" -- 5590
           ,x"0887" -- 5592
           ,x"15cc" -- 5594
           ,x"06a0" -- 5596
           ,x"bf34" -- 5598
           ,x"0587" -- 559A
           ,x"16fc" -- 559C
           ,x"d008" -- 559E
           ,x"0240" -- 55A0
           ,x"80ff" -- 55A2
           ,x"b004" -- 55A4
           ,x"0380" -- 55A6
           ,x"9838" -- 55A8
           ,x"ad1f" -- 55AA
           ,x"1616" -- 55AC
           ,x"0420" -- 55AE
           ,x"b540" -- 55B0
           ,x"0280" -- 55B2
           ,x"3f00" -- 55B4
           ,x"1611" -- 55B6
           ,x"06a0" -- 55B8
           ,x"c1b0" -- 55BA
           ,x"c041" -- 55BC
           ,x"1501" -- 55BE
           ,x"04c1" -- 55C0
           ,x"c001" -- 55C2
           ,x"0931" -- 55C4
           ,x"a081" -- 55C6
           ,x"0201" -- 55C8
           ,x"8000" -- 55CA
           ,x"0b01" -- 55CC
           ,x"4481" -- 55CE
           ,x"c0c3" -- 55D0
           ,x"1301" -- 55D2
           ,x"e481" -- 55D4
           ,x"0460" -- 55D6
           ,x"aefc" -- 55D8
           ,x"0460" -- 55DA
           ,x"97b2" -- 55DC
           ,x"c041" -- 55DE
           ,x"1501" -- 55E0
           ,x"04c1" -- 55E2
           ,x"c001" -- 55E4
           ,x"0931" -- 55E6
           ,x"a081" -- 55E8
           ,x"0201" -- 55EA
           ,x"8000" -- 55EC
           ,x"0b01" -- 55EE
           ,x"c092" -- 55F0
           ,x"2081" -- 55F2
           ,x"1602" -- 55F4
           ,x"05a0" -- 55F6
           ,x"ef6a" -- 55F8
           ,x"0460" -- 55FA
           ,x"b6be" -- 55FC
           ,x"c3a0" -- 55FE
           ,x"ede4" -- 5600
           ,x"1634" -- 5602
           ,x"c1e0" -- 5604
           ,x"ed04" -- 5606
           ,x"0420" -- 5608
           ,x"b284" -- 560A
           ,x"1000" -- 560C
           ,x"100b" -- 560E
           ,x"06a0" -- 5610
           ,x"a2a6" -- 5612
           ,x"c1e0" -- 5614
           ,x"ed04" -- 5616
           ,x"0720" -- 5618
           ,x"ede2" -- 561A
           ,x"06a0" -- 561C
           ,x"ac2c" -- 561E
           ,x"0420" -- 5620
           ,x"8170" -- 5622
           ,x"101b" -- 5624
           ,x"0420" -- 5626
           ,x"8d70" -- 5628
           ,x"000d" -- 562A
           ,x"c80b" -- 562C
           ,x"edd0" -- 562E
           ,x"0206" -- 5630
           ,x"0064" -- 5632
           ,x"c1e0" -- 5634
           ,x"ed04" -- 5636
           ,x"c0c7" -- 5638
           ,x"c046" -- 563A
           ,x"04f3" -- 563C
           ,x"0641" -- 563E
           ,x"15fd" -- 5640
           ,x"c060" -- 5642
           ,x"ede0" -- 5644
           ,x"1311" -- 5646
           ,x"a060" -- 5648
           ,x"edee" -- 564A
           ,x"1131" -- 564C
           ,x"c820" -- 564E
           ,x"801a" -- 5650
           ,x"ef9e" -- 5652
           ,x"0420" -- 5654
           ,x"b05a" -- 5656
           ,x"dde0" -- 5658
           ,x"c0e4" -- 565A
           ,x"0420" -- 565C
           ,x"8174" -- 565E
           ,x"0206" -- 5660
           ,x"0064" -- 5662
           ,x"a1a0" -- 5664
           ,x"ed04" -- 5666
           ,x"6187" -- 5668
           ,x"04cf" -- 566A
           ,x"0420" -- 566C
           ,x"8198" -- 566E
           ,x"0280" -- 5670
           ,x"2000" -- 5672
           ,x"1401" -- 5674
           ,x"04cf" -- 5676
           ,x"06a0" -- 5678
           ,x"872c" -- 567A
           ,x"5a17" -- 567C
           ,x"c105" -- 567E
           ,x"3909" -- 5680
           ,x"2308" -- 5682
           ,x"7016" -- 5684
           ,x"170c" -- 5686
           ,x"f80a" -- 5688
           ,x"1a0d" -- 568A
           ,x"287f" -- 568C
           ,x"0000" -- 568E
           ,x"0280" -- 5690
           ,x"2000" -- 5692
           ,x"1a09" -- 5694
           ,x"d157" -- 5696
           ,x"1602" -- 5698
           ,x"0606" -- 569A
           ,x"1104" -- 569C
           ,x"c3cf" -- 569E
           ,x"165f" -- 56A0
           ,x"ddc0" -- 56A2
           ,x"1002" -- 56A4
           ,x"0586" -- 56A6
           ,x"10e1" -- 56A8
           ,x"0420" -- 56AA
           ,x"816c" -- 56AC
           ,x"10de" -- 56AE
           ,x"ddd7" -- 56B0
           ,x"1304" -- 56B2
           ,x"0420" -- 56B4
           ,x"818c" -- 56B6
           ,x"0900" -- 56B8
           ,x"10fa" -- 56BA
           ,x"c2e0" -- 56BC
           ,x"edd0" -- 56BE
           ,x"045b" -- 56C0
           ,x"81e0" -- 56C2
           ,x"ed04" -- 56C4
           ,x"13f0" -- 56C6
           ,x"0607" -- 56C8
           ,x"100d" -- 56CA
           ,x"04cf" -- 56CC
           ,x"81e0" -- 56CE
           ,x"ed04" -- 56D0
           ,x"13ea" -- 56D2
           ,x"0607" -- 56D4
           ,x"d5e0" -- 56D6
           ,x"c0e4" -- 56D8
           ,x"0420" -- 56DA
           ,x"818c" -- 56DC
           ,x"0800" -- 56DE
           ,x"0420" -- 56E0
           ,x"818c" -- 56E2
           ,x"2000" -- 56E4
           ,x"0420" -- 56E6
           ,x"818c" -- 56E8
           ,x"0800" -- 56EA
           ,x"10bf" -- 56EC
           ,x"d037" -- 56EE
           ,x"16dc" -- 56F0
           ,x"0607" -- 56F2
           ,x"10d9" -- 56F4
           ,x"c0e0" -- 56F6
           ,x"804a" -- 56F8
           ,x"1302" -- 56FA
           ,x"0460" -- 56FC
           ,x"8124" -- 56FE
           ,x"c0db" -- 5700
           ,x"0607" -- 5702
           ,x"c147" -- 5704
           ,x"06a0" -- 5706
           ,x"8d0a" -- 5708
           ,x"c1a0" -- 570A
           ,x"ed02" -- 570C
           ,x"0420" -- 570E
           ,x"8170" -- 5710
           ,x"0420" -- 5712
           ,x"8174" -- 5714
           ,x"0420" -- 5716
           ,x"818c" -- 5718
           ,x"0d00" -- 571A
           ,x"c1e0" -- 571C
           ,x"ed04" -- 571E
           ,x"04cf" -- 5720
           ,x"8147" -- 5722
           ,x"14a3" -- 5724
           ,x"04c0" -- 5726
           ,x"d037" -- 5728
           ,x"0420" -- 572A
           ,x"816c" -- 572C
           ,x"10f9" -- 572E
           ,x"d5d7" -- 5730
           ,x"13ba" -- 5732
           ,x"c047" -- 5734
           ,x"dde7" -- 5736
           ,x"0001" -- 5738
           ,x"16fd" -- 573A
           ,x"d451" -- 573C
           ,x"1302" -- 573E
           ,x"0420" -- 5740
           ,x"8178" -- 5742
           ,x"0420" -- 5744
           ,x"818c" -- 5746
           ,x"2000" -- 5748
           ,x"61c1" -- 574A
           ,x"0420" -- 574C
           ,x"818c" -- 574E
           ,x"0800" -- 5750
           ,x"0607" -- 5752
           ,x"16fb" -- 5754
           ,x"c1c1" -- 5756
           ,x"0586" -- 5758
           ,x"1088" -- 575A
           ,x"070f" -- 575C
           ,x"1086" -- 575E
           ,x"0606" -- 5760
           ,x"11a1" -- 5762
           ,x"13a0" -- 5764
           ,x"c047" -- 5766
           ,x"ddd7" -- 5768
           ,x"16fe" -- 576A
           ,x"d5e7" -- 576C
           ,x"ffff" -- 576E
           ,x"0607" -- 5770
           ,x"8047" -- 5772
           ,x"1bfb" -- 5774
           ,x"ddc0" -- 5776
           ,x"0420" -- 5778
           ,x"8178" -- 577A
           ,x"0581" -- 577C
           ,x"d031" -- 577E
           ,x"13ec" -- 5780
           ,x"0420" -- 5782
           ,x"818c" -- 5784
           ,x"0800" -- 5786
           ,x"10fa" -- 5788
           ,x"0202" -- 578A
           ,x"c1a2" -- 578C
           ,x"0812" -- 578E
           ,x"a083" -- 5790
           ,x"0a12" -- 5792
           ,x"c812" -- 5794
           ,x"edf8" -- 5796
           ,x"c820" -- 5798
           ,x"800a" -- 579A
           ,x"ef7e" -- 579C
           ,x"0420" -- 579E
           ,x"bd84" -- 57A0
           ,x"045b" -- 57A2
           ,x"4120" -- 57A4
           ,x"4140" -- 57A6
           ,x"4180" -- 57A8
           ,x"9838" -- 57AA
           ,x"ad1f" -- 57AC
           ,x"1611" -- 57AE
           ,x"c820" -- 57B0
           ,x"801a" -- 57B2
           ,x"ef9e" -- 57B4
           ,x"0420" -- 57B6
           ,x"b558" -- 57B8
           ,x"0280" -- 57BA
           ,x"4b00" -- 57BC
           ,x"1609" -- 57BE
           ,x"9e20" -- 57C0
           ,x"ab26" -- 57C2
           ,x"1608" -- 57C4
           ,x"c820" -- 57C6
           ,x"801e" -- 57C8
           ,x"ef9e" -- 57CA
           ,x"0420" -- 57CC
           ,x"b558" -- 57CE
           ,x"045b" -- 57D0
           ,x"0460" -- 57D2
           ,x"97b2" -- 57D4
           ,x"0460" -- 57D6
           ,x"9802" -- 57D8
           ,x"0420" -- 57DA
           ,x"8d70" -- 57DC
           ,x"001a" -- 57DE
           ,x"c28b" -- 57E0
           ,x"06a0" -- 57E2
           ,x"c4d0" -- 57E4
           ,x"10f9" -- 57E6
           ,x"c0c3" -- 57E8
           ,x"16f7" -- 57EA
           ,x"d820" -- 57EC
           ,x"c8e0" -- 57EE
           ,x"ef68" -- 57F0
           ,x"0961" -- 57F2
           ,x"0221" -- 57F4
           ,x"ff00" -- 57F6
           ,x"c092" -- 57F8
           ,x"0200" -- 57FA
           ,x"0080" -- 57FC
           ,x"2080" -- 57FE
           ,x"1308" -- 5800
           ,x"04c3" -- 5802
           ,x"0583" -- 5804
           ,x"0910" -- 5806
           ,x"2080" -- 5808
           ,x"16fc" -- 580A
           ,x"6043" -- 580C
           ,x"06a0" -- 580E
           ,x"c18a" -- 5810
           ,x"c081" -- 5812
           ,x"c820" -- 5814
           ,x"8012" -- 5816
           ,x"ef7e" -- 5818
           ,x"0420" -- 581A
           ,x"bc32" -- 581C
           ,x"c820" -- 581E
           ,x"c2ec" -- 5820
           ,x"ef7e" -- 5822
           ,x"0420" -- 5824
           ,x"bc4e" -- 5826
           ,x"0200" -- 5828
           ,x"c2fe" -- 582A
           ,x"c060" -- 582C
           ,x"ef68" -- 582E
           ,x"1504" -- 5830
           ,x"1303" -- 5832
           ,x"0200" -- 5834
           ,x"c2f6" -- 5836
           ,x"0602" -- 5838
           ,x"c820" -- 583A
           ,x"8012" -- 583C
           ,x"ef7e" -- 583E
           ,x"0420" -- 5840
           ,x"bc3e" -- 5842
           ,x"c800" -- 5844
           ,x"ef7e" -- 5846
           ,x"0420" -- 5848
           ,x"bc4a" -- 584A
           ,x"c820" -- 584C
           ,x"8000" -- 584E
           ,x"ef7e" -- 5850
           ,x"0420" -- 5852
           ,x"bc32" -- 5854
           ,x"c820" -- 5856
           ,x"8012" -- 5858
           ,x"ef7e" -- 585A
           ,x"0420" -- 585C
           ,x"bc3e" -- 585E
           ,x"c800" -- 5860
           ,x"ef7e" -- 5862
           ,x"0420" -- 5864
           ,x"bc4e" -- 5866
           ,x"c820" -- 5868
           ,x"8000" -- 586A
           ,x"ef7e" -- 586C
           ,x"0420" -- 586E
           ,x"beac" -- 5870
           ,x"c820" -- 5872
           ,x"8000" -- 5874
           ,x"ef7e" -- 5876
           ,x"0420" -- 5878
           ,x"bc32" -- 587A
           ,x"06a0" -- 587C
           ,x"c4f4" -- 587E
           ,x"c2fc" -- 5880
           ,x"c820" -- 5882
           ,x"8002" -- 5884
           ,x"ef7e" -- 5886
           ,x"0420" -- 5888
           ,x"bc32" -- 588A
           ,x"06a0" -- 588C
           ,x"c512" -- 588E
           ,x"c316" -- 5890
           ,x"c820" -- 5892
           ,x"8002" -- 5894
           ,x"ef7e" -- 5896
           ,x"0420" -- 5898
           ,x"beac" -- 589A
           ,x"c820" -- 589C
           ,x"8000" -- 589E
           ,x"ef7e" -- 58A0
           ,x"0420" -- 58A2
           ,x"bd84" -- 58A4
           ,x"c820" -- 58A6
           ,x"8012" -- 58A8
           ,x"ef7e" -- 58AA
           ,x"0420" -- 58AC
           ,x"bc32" -- 58AE
           ,x"0200" -- 58B0
           ,x"8c00" -- 58B2
           ,x"c082" -- 58B4
           ,x"1102" -- 58B6
           ,x"0910" -- 58B8
           ,x"1002" -- 58BA
           ,x"0502" -- 58BC
           ,x"0810" -- 58BE
           ,x"c042" -- 58C0
           ,x"04c2" -- 58C2
           ,x"c820" -- 58C4
           ,x"8016" -- 58C6
           ,x"ef7e" -- 58C8
           ,x"0420" -- 58CA
           ,x"bc3e" -- 58CC
           ,x"0420" -- 58CE
           ,x"bd46" -- 58D0
           ,x"c820" -- 58D2
           ,x"c2ee" -- 58D4
           ,x"ef7e" -- 58D6
           ,x"0420" -- 58D8
           ,x"bd84" -- 58DA
           ,x"c820" -- 58DC
           ,x"8012" -- 58DE
           ,x"ef7e" -- 58E0
           ,x"0420" -- 58E2
           ,x"bc4a" -- 58E4
           ,x"0202" -- 58E6
           ,x"ef68" -- 58E8
           ,x"045a" -- 58EA
           ,x"c2f0" -- 58EC
           ,x"c32a" -- 58EE
           ,x"40b5" -- 58F0
           ,x"04f3" -- 58F2
           ,x"33fa" -- 58F4
           ,x"4080" -- 58F6
           ,x"0000" -- 58F8
           ,x"0000" -- 58FA
           ,x"0003" -- 58FC
           ,x"4110" -- 58FE
           ,x"0000" -- 5900
           ,x"0000" -- 5902
           ,x"c214" -- 5904
           ,x"bbc5" -- 5906
           ,x"dcdb" -- 5908
           ,x"423d" -- 590A
           ,x"c2d5" -- 590C
           ,x"31f0" -- 590E
           ,x"c22d" -- 5910
           ,x"165c" -- 5912
           ,x"4be0" -- 5914
           ,x"0002" -- 5916
           ,x"c212" -- 5918
           ,x"53ef" -- 591A
           ,x"500e" -- 591C
           ,x"425d" -- 591E
           ,x"76c2" -- 5920
           ,x"314a" -- 5922
           ,x"c25a" -- 5924
           ,x"2cb8" -- 5926
           ,x"97bf" -- 5928
           ,x"40b1" -- 592A
           ,x"7217" -- 592C
           ,x"f7d2" -- 592E
           ,x"070d" -- 5930
           ,x"1001" -- 5932
           ,x"04cd" -- 5934
           ,x"0420" -- 5936
           ,x"81a8" -- 5938
           ,x"06a0" -- 593A
           ,x"8724" -- 593C
           ,x"1838" -- 593E
           ,x"1600" -- 5940
           ,x"163c" -- 5942
           ,x"1647" -- 5944
           ,x"0000" -- 5946
           ,x"0608" -- 5948
           ,x"06a0" -- 594A
           ,x"c390" -- 594C
           ,x"d80f" -- 594E
           ,x"ef42" -- 5950
           ,x"d80e" -- 5952
           ,x"ef43" -- 5954
           ,x"0280" -- 5956
           ,x"3800" -- 5958
           ,x"1309" -- 595A
           ,x"c34d" -- 595C
           ,x"1303" -- 595E
           ,x"0420" -- 5960
           ,x"8c68" -- 5962
           ,x"1002" -- 5964
           ,x"0420" -- 5966
           ,x"8c72" -- 5968
           ,x"0460" -- 596A
           ,x"aefc" -- 596C
           ,x"06a0" -- 596E
           ,x"c390" -- 5970
           ,x"d80f" -- 5972
           ,x"ed92" -- 5974
           ,x"d80e" -- 5976
           ,x"ed93" -- 5978
           ,x"c34d" -- 597A
           ,x"1606" -- 597C
           ,x"0420" -- 597E
           ,x"c3be" -- 5980
           ,x"0280" -- 5982
           ,x"3800" -- 5984
           ,x"13f3" -- 5986
           ,x"10f0" -- 5988
           ,x"0420" -- 598A
           ,x"c3b4" -- 598C
           ,x"10f9" -- 598E
           ,x"c820" -- 5990
           ,x"802a" -- 5992
           ,x"ef9e" -- 5994
           ,x"0420" -- 5996
           ,x"b558" -- 5998
           ,x"06cf" -- 599A
           ,x"0280" -- 599C
           ,x"3f00" -- 599E
           ,x"1607" -- 59A0
           ,x"c820" -- 59A2
           ,x"8028" -- 59A4
           ,x"ef9e" -- 59A6
           ,x"0420" -- 59A8
           ,x"b558" -- 59AA
           ,x"06ce" -- 59AC
           ,x"045b" -- 59AE
           ,x"0460" -- 59B0
           ,x"aef2" -- 59B2
           ,x"ef20" -- 59B4
           ,x"c3b8" -- 59B6
           ,x"0200" -- 59B8
           ,x"8c68" -- 59BA
           ,x"1004" -- 59BC
           ,x"ef20" -- 59BE
           ,x"c3c2" -- 59C0
           ,x"0200" -- 59C2
           ,x"8c72" -- 59C4
           ,x"070b" -- 59C6
           ,x"070a" -- 59C8
           ,x"0709" -- 59CA
           ,x"04c3" -- 59CC
           ,x"04c4" -- 59CE
           ,x"d820" -- 59D0
           ,x"ef42" -- 59D2
           ,x"ef29" -- 59D4
           ,x"d820" -- 59D6
           ,x"ed92" -- 59D8
           ,x"ef27" -- 59DA
           ,x"6103" -- 59DC
           ,x"0744" -- 59DE
           ,x"1101" -- 59E0
           ,x"050a" -- 59E2
           ,x"d820" -- 59E4
           ,x"ef43" -- 59E6
           ,x"ef27" -- 59E8
           ,x"04c5" -- 59EA
           ,x"d820" -- 59EC
           ,x"ed93" -- 59EE
           ,x"ef2b" -- 59F0
           ,x"60c5" -- 59F2
           ,x"0743" -- 59F4
           ,x"1101" -- 59F6
           ,x"0509" -- 59F8
           ,x"80c4" -- 59FA
           ,x"1508" -- 59FC
           ,x"2903" -- 59FE
           ,x"28c4" -- 5A00
           ,x"2903" -- 5A02
           ,x"d160" -- 5A04
           ,x"ed93" -- 5A06
           ,x"d1a0" -- 5A08
           ,x"ed92" -- 5A0A
           ,x"1008" -- 5A0C
           ,x"d160" -- 5A0E
           ,x"ed92" -- 5A10
           ,x"d1a0" -- 5A12
           ,x"ed93" -- 5A14
           ,x"2a89" -- 5A16
           ,x"2a4a" -- 5A18
           ,x"2a89" -- 5A1A
           ,x"05cb" -- 5A1C
           ,x"0985" -- 5A1E
           ,x"0986" -- 5A20
           ,x"0a53" -- 5A22
           ,x"04c2" -- 5A24
           ,x"3c84" -- 5A26
           ,x"c1c2" -- 5A28
           ,x"c083" -- 5A2A
           ,x"04c3" -- 5A2C
           ,x"1901" -- 5A2E
           ,x"1003" -- 5A30
           ,x"3c84" -- 5A32
           ,x"c0c2" -- 5A34
           ,x"c087" -- 5A36
           ,x"0207" -- 5A38
           ,x"0010" -- 5A3A
           ,x"04c8" -- 5A3C
           ,x"04cc" -- 5A3E
           ,x"810c" -- 5A40
           ,x"1b1d" -- 5A42
           ,x"058c" -- 5A44
           ,x"c2cb" -- 5A46
           ,x"1107" -- 5A48
           ,x"d820" -- 5A4A
           ,x"ef2b" -- 5A4C
           ,x"ef42" -- 5A4E
           ,x"d820" -- 5A50
           ,x"ef2d" -- 5A52
           ,x"ef43" -- 5A54
           ,x"1006" -- 5A56
           ,x"d820" -- 5A58
           ,x"ef2d" -- 5A5A
           ,x"ef42" -- 5A5C
           ,x"d820" -- 5A5E
           ,x"ef2b" -- 5A60
           ,x"ef43" -- 5A62
           ,x"0410" -- 5A64
           ,x"a203" -- 5A66
           ,x"1701" -- 5A68
           ,x"0587" -- 5A6A
           ,x"a1c2" -- 5A6C
           ,x"0287" -- 5A6E
           ,x"0020" -- 5A70
           ,x"1a03" -- 5A72
           ,x"0227" -- 5A74
           ,x"ffe0" -- 5A76
           ,x"a18a" -- 5A78
           ,x"a149" -- 5A7A
           ,x"10e1" -- 5A7C
           ,x"d820" -- 5A7E
           ,x"ed92" -- 5A80
           ,x"ef42" -- 5A82
           ,x"d820" -- 5A84
           ,x"ed93" -- 5A86
           ,x"ef43" -- 5A88
           ,x"0380" -- 5A8A
           ,x"c060" -- 5A8C
           ,x"ef68" -- 5A8E
           ,x"a041" -- 5A90
           ,x"0281" -- 5A92
           ,x"8900" -- 5A94
           ,x"1b1a" -- 5A96
           ,x"c820" -- 5A98
           ,x"8012" -- 5A9A
           ,x"ef7e" -- 5A9C
           ,x"0420" -- 5A9E
           ,x"bc32" -- 5AA0
           ,x"c820" -- 5AA2
           ,x"c83a" -- 5AA4
           ,x"ef7e" -- 5AA6
           ,x"0420" -- 5AA8
           ,x"bf7c" -- 5AAA
           ,x"c060" -- 5AAC
           ,x"ef6c" -- 5AAE
           ,x"c0a0" -- 5AB0
           ,x"ef68" -- 5AB2
           ,x"1501" -- 5AB4
           ,x"0501" -- 5AB6
           ,x"0420" -- 5AB8
           ,x"bd46" -- 5ABA
           ,x"0420" -- 5ABC
           ,x"bd0c" -- 5ABE
           ,x"c820" -- 5AC0
           ,x"8012" -- 5AC2
           ,x"ef7e" -- 5AC4
           ,x"0420" -- 5AC6
           ,x"bc4a" -- 5AC8
           ,x"045b" -- 5ACA
           ,x"0460" -- 5ACC
           ,x"bc10" -- 5ACE
           ,x"c802" -- 5AD0
           ,x"ef7e" -- 5AD2
           ,x"0420" -- 5AD4
           ,x"bc3e" -- 5AD6
           ,x"0420" -- 5AD8
           ,x"bd1a" -- 5ADA
           ,x"0202" -- 5ADC
           ,x"ef68" -- 5ADE
           ,x"c0d2" -- 5AE0
           ,x"1307" -- 5AE2
           ,x"09f3" -- 5AE4
           ,x"1302" -- 5AE6
           ,x"0420" -- 5AE8
           ,x"bd0c" -- 5AEA
           ,x"05cb" -- 5AEC
           ,x"04c1" -- 5AEE
           ,x"d052" -- 5AF0
           ,x"045b" -- 5AF2
           ,x"c820" -- 5AF4
           ,x"8012" -- 5AF6
           ,x"ef7e" -- 5AF8
           ,x"0420" -- 5AFA
           ,x"bc32" -- 5AFC
           ,x"c820" -- 5AFE
           ,x"8012" -- 5B00
           ,x"ef7e" -- 5B02
           ,x"0420" -- 5B04
           ,x"bd84" -- 5B06
           ,x"c820" -- 5B08
           ,x"8012" -- 5B0A
           ,x"ef7e" -- 5B0C
           ,x"0420" -- 5B0E
           ,x"bc32" -- 5B10
           ,x"c03b" -- 5B12
           ,x"c070" -- 5B14
           ,x"c800" -- 5B16
           ,x"ef7e" -- 5B18
           ,x"0420" -- 5B1A
           ,x"bc3e" -- 5B1C
           ,x"c820" -- 5B1E
           ,x"8012" -- 5B20
           ,x"ef7e" -- 5B22
           ,x"0420" -- 5B24
           ,x"bd84" -- 5B26
           ,x"0220" -- 5B28
           ,x"0006" -- 5B2A
           ,x"c800" -- 5B2C
           ,x"ef7e" -- 5B2E
           ,x"0420" -- 5B30
           ,x"bc4a" -- 5B32
           ,x"0601" -- 5B34
           ,x"16f3" -- 5B36
           ,x"045b" -- 5B38
           ,x"c101" -- 5B3A
           ,x"c800" -- 5B3C
           ,x"ef66" -- 5B3E
           ,x"06a0" -- 5B40
           ,x"c1e0" -- 5B42
           ,x"c820" -- 5B44
           ,x"8012" -- 5B46
           ,x"ef7e" -- 5B48
           ,x"0420" -- 5B4A
           ,x"bc32" -- 5B4C
           ,x"c804" -- 5B4E
           ,x"ef7e" -- 5B50
           ,x"0420" -- 5B52
           ,x"bc3e" -- 5B54
           ,x"0420" -- 5B56
           ,x"bd1a" -- 5B58
           ,x"c820" -- 5B5A
           ,x"8012" -- 5B5C
           ,x"ef7e" -- 5B5E
           ,x"0420" -- 5B60
           ,x"bd84" -- 5B62
           ,x"06a0" -- 5B64
           ,x"baaa" -- 5B66
           ,x"c020" -- 5B68
           ,x"ef66" -- 5B6A
           ,x"0460" -- 5B6C
           ,x"b82e" -- 5B6E
           ,x"c020" -- 5B70
           ,x"ed00" -- 5B72
           ,x"c0c0" -- 5B74
           ,x"0ab3" -- 5B76
           ,x"a0c0" -- 5B78
           ,x"0a23" -- 5B7A
           ,x"a003" -- 5B7C
           ,x"0220" -- 5B7E
           ,x"3619" -- 5B80
           ,x"c800" -- 5B82
           ,x"ed00" -- 5B84
           ,x"045b" -- 5B86
           ,x"ef68" -- 5B88
           ,x"c58c" -- 5B8A
           ,x"06a0" -- 5B8C
           ,x"c570" -- 5B8E
           ,x"c040" -- 5B90
           ,x"06a0" -- 5B92
           ,x"c570" -- 5B94
           ,x"c080" -- 5B96
           ,x"0200" -- 5B98
           ,x"4200" -- 5B9A
           ,x"0460" -- 5B9C
           ,x"bd4a" -- 5B9E
           ,x"c28b" -- 5BA0
           ,x"06a0" -- 5BA2
           ,x"c4d0" -- 5BA4
           ,x"1003" -- 5BA6
           ,x"0203" -- 5BA8
           ,x"0001" -- 5BAA
           ,x"100b" -- 5BAC
           ,x"c820" -- 5BAE
           ,x"c63a" -- 5BB0
           ,x"ef7e" -- 5BB2
           ,x"0420" -- 5BB4
           ,x"bc3e" -- 5BB6
           ,x"103c" -- 5BB8
           ,x"c28b" -- 5BBA
           ,x"06a0" -- 5BBC
           ,x"c4d0" -- 5BBE
           ,x"1038" -- 5BC0
           ,x"0a13" -- 5BC2
           ,x"c820" -- 5BC4
           ,x"c638" -- 5BC6
           ,x"ef7e" -- 5BC8
           ,x"0420" -- 5BCA
           ,x"bd84" -- 5BCC
           ,x"06a0" -- 5BCE
           ,x"c48c" -- 5BD0
           ,x"a043" -- 5BD2
           ,x"0911" -- 5BD4
           ,x"170f" -- 5BD6
           ,x"c820" -- 5BD8
           ,x"8012" -- 5BDA
           ,x"ef7e" -- 5BDC
           ,x"0420" -- 5BDE
           ,x"bc32" -- 5BE0
           ,x"c820" -- 5BE2
           ,x"c63a" -- 5BE4
           ,x"ef7e" -- 5BE6
           ,x"0420" -- 5BE8
           ,x"bc3e" -- 5BEA
           ,x"c820" -- 5BEC
           ,x"8012" -- 5BEE
           ,x"ef7e" -- 5BF0
           ,x"0420" -- 5BF2
           ,x"bc4e" -- 5BF4
           ,x"0911" -- 5BF6
           ,x"1702" -- 5BF8
           ,x"0420" -- 5BFA
           ,x"bd0c" -- 5BFC
           ,x"c820" -- 5BFE
           ,x"8000" -- 5C00
           ,x"ef7e" -- 5C02
           ,x"0420" -- 5C04
           ,x"bc32" -- 5C06
           ,x"06a0" -- 5C08
           ,x"c4f4" -- 5C0A
           ,x"c642" -- 5C0C
           ,x"c820" -- 5C0E
           ,x"8002" -- 5C10
           ,x"ef7e" -- 5C12
           ,x"0420" -- 5C14
           ,x"bc32" -- 5C16
           ,x"06a0" -- 5C18
           ,x"c512" -- 5C1A
           ,x"c656" -- 5C1C
           ,x"c820" -- 5C1E
           ,x"8002" -- 5C20
           ,x"ef7e" -- 5C22
           ,x"0420" -- 5C24
           ,x"beac" -- 5C26
           ,x"c820" -- 5C28
           ,x"8000" -- 5C2A
           ,x"ef7e" -- 5C2C
           ,x"0420" -- 5C2E
           ,x"bd84" -- 5C30
           ,x"0202" -- 5C32
           ,x"ef68" -- 5C34
           ,x"045a" -- 5C36
           ,x"c63c" -- 5C38
           ,x"c644" -- 5C3A
           ,x"40a2" -- 5C3C
           ,x"f983" -- 5C3E
           ,x"6e4e" -- 5C40
           ,x"0002" -- 5C42
           ,x"4110" -- 5C44
           ,x"0000" -- 5C46
           ,x"0000" -- 5C48
           ,x"4273" -- 5C4A
           ,x"4dca" -- 5C4C
           ,x"815d" -- 5C4E
           ,x"4411" -- 5C50
           ,x"7825" -- 5C52
           ,x"55b4" -- 5C54
           ,x"0005" -- 5C56
           ,x"be95" -- 5C58
           ,x"3606" -- 5C5A
           ,x"2dee" -- 5C5C
           ,x"4041" -- 5C5E
           ,x"e3f5" -- 5C60
           ,x"31b8" -- 5C62
           ,x"c1c6" -- 5C64
           ,x"5036" -- 5C66
           ,x"51d0" -- 5C68
           ,x"4311" -- 5C6A
           ,x"b7c5" -- 5C6C
           ,x"5a8f" -- 5C6E
           ,x"c3a9" -- 5C70
           ,x"3ba0" -- 5C72
           ,x"c828" -- 5C74
           ,x"441b" -- 5C76
           ,x"70d4" -- 5C78
           ,x"8bb5" -- 5C7A
           ,x"06a0" -- 5C7C
           ,x"c4d0" -- 5C7E
           ,x"103d" -- 5C80
           ,x"c0c3" -- 5C82
           ,x"1641" -- 5C84
           ,x"c820" -- 5C86
           ,x"8000" -- 5C88
           ,x"ef7e" -- 5C8A
           ,x"0420" -- 5C8C
           ,x"bc32" -- 5C8E
           ,x"0200" -- 5C90
           ,x"4000" -- 5C92
           ,x"6040" -- 5C94
           ,x"d800" -- 5C96
           ,x"ef68" -- 5C98
           ,x"c820" -- 5C9A
           ,x"c70e" -- 5C9C
           ,x"ef7e" -- 5C9E
           ,x"0420" -- 5CA0
           ,x"bd84" -- 5CA2
           ,x"c820" -- 5CA4
           ,x"c710" -- 5CA6
           ,x"ef7e" -- 5CA8
           ,x"0420" -- 5CAA
           ,x"bc4a" -- 5CAC
           ,x"0991" -- 5CAE
           ,x"1705" -- 5CB0
           ,x"c820" -- 5CB2
           ,x"c714" -- 5CB4
           ,x"ef7e" -- 5CB6
           ,x"0420" -- 5CB8
           ,x"bd84" -- 5CBA
           ,x"06c1" -- 5CBC
           ,x"b801" -- 5CBE
           ,x"ef68" -- 5CC0
           ,x"0201" -- 5CC2
           ,x"0004" -- 5CC4
           ,x"c820" -- 5CC6
           ,x"8012" -- 5CC8
           ,x"ef7e" -- 5CCA
           ,x"0420" -- 5CCC
           ,x"bc32" -- 5CCE
           ,x"c820" -- 5CD0
           ,x"8000" -- 5CD2
           ,x"ef7e" -- 5CD4
           ,x"0420" -- 5CD6
           ,x"bc3e" -- 5CD8
           ,x"c820" -- 5CDA
           ,x"8012" -- 5CDC
           ,x"ef7e" -- 5CDE
           ,x"0420" -- 5CE0
           ,x"beac" -- 5CE2
           ,x"c820" -- 5CE4
           ,x"8012" -- 5CE6
           ,x"ef7e" -- 5CE8
           ,x"0420" -- 5CEA
           ,x"bc4a" -- 5CEC
           ,x"c820" -- 5CEE
           ,x"c712" -- 5CF0
           ,x"ef7e" -- 5CF2
           ,x"0420" -- 5CF4
           ,x"bd84" -- 5CF6
           ,x"0601" -- 5CF8
           ,x"16e5" -- 5CFA
           ,x"0202" -- 5CFC
           ,x"ef68" -- 5CFE
           ,x"44a0" -- 5D00
           ,x"bfca" -- 5D02
           ,x"06a0" -- 5D04
           ,x"b6ac" -- 5D06
           ,x"0420" -- 5D08
           ,x"8d70" -- 5D0A
           ,x"0019" -- 5D0C
           ,x"c716" -- 5D0E
           ,x"c71c" -- 5D10
           ,x"c722" -- 5D12
           ,x"c728" -- 5D14
           ,x"40e4" -- 5D16
           ,x"f92a" -- 5D18
           ,x"f9a8" -- 5D1A
           ,x"4039" -- 5D1C
           ,x"3e4e" -- 5D1E
           ,x"f028" -- 5D20
           ,x"4080" -- 5D22
           ,x"0000" -- 5D24
           ,x"0000" -- 5D26
           ,x"4140" -- 5D28
           ,x"0000" -- 5D2A
           ,x"0000" -- 5D2C
           ,x"06a0" -- 5D2E
           ,x"a364" -- 5D30
           ,x"0202" -- 5D32
           ,x"c75c" -- 5D34
           ,x"c288" -- 5D36
           ,x"c0f2" -- 5D38
           ,x"130d" -- 5D3A
           ,x"c132" -- 5D3C
           ,x"d038" -- 5D3E
           ,x"1305" -- 5D40
           ,x"9032" -- 5D42
           ,x"13fc" -- 5D44
           ,x"c083" -- 5D46
           ,x"c20a" -- 5D48
           ,x"10f6" -- 5D4A
           ,x"d012" -- 5D4C
           ,x"16fb" -- 5D4E
           ,x"2fa0" -- 5D50
           ,x"c8b9" -- 5D52
           ,x"0454" -- 5D54
           ,x"0420" -- 5D56
           ,x"8d70" -- 5D58
           ,x"0029" -- 5D5A
           ,x"c764" -- 5D5C
           ,x"c786" -- 5D5E
           ,x"4449" -- 5D60
           ,x"5200" -- 5D62
           ,x"c76e" -- 5D64
           ,x"c78e" -- 5D66
           ,x"5341" -- 5D68
           ,x"5645" -- 5D6A
           ,x"0000" -- 5D6C
           ,x"c778" -- 5D6E
           ,x"c7e2" -- 5D70
           ,x"4c4f" -- 5D72
           ,x"4144" -- 5D74
           ,x"0000" -- 5D76
           ,x"c784" -- 5D78
           ,x"c830" -- 5D7A
           ,x"4445" -- 5D7C
           ,x"4c45" -- 5D7E
           ,x"5445" -- 5D80
           ,x"0000" -- 5D82
           ,x"0000" -- 5D84
           ,x"0420" -- 5D86
           ,x"1562" -- 5D88
           ,x"0460" -- 5D8A
           ,x"8116" -- 5D8C
           ,x"c060" -- 5D8E
           ,x"ed0e" -- 5D90
           ,x"c241" -- 5D92
           ,x"0221" -- 5D94
           ,x"fff8" -- 5D96
           ,x"c460" -- 5D98
           ,x"edd2" -- 5D9A
           ,x"6c49" -- 5D9C
           ,x"c460" -- 5D9E
           ,x"edd4" -- 5DA0
           ,x"6c49" -- 5DA2
           ,x"c460" -- 5DA4
           ,x"edd8" -- 5DA6
           ,x"6c60" -- 5DA8
           ,x"edd6" -- 5DAA
           ,x"c460" -- 5DAC
           ,x"edd8" -- 5DAE
           ,x"6449" -- 5DB0
           ,x"0207" -- 5DB2
           ,x"000a" -- 5DB4
           ,x"a447" -- 5DB6
           ,x"0229" -- 5DB8
           ,x"fff6" -- 5DBA
           ,x"c660" -- 5DBC
           ,x"c840" -- 5DBE
           ,x"0420" -- 5DC0
           ,x"8184" -- 5DC2
           ,x"c8c1" -- 5DC4
           ,x"06a0" -- 5DC6
           ,x"8754" -- 5DC8
           ,x"10fa" -- 5DCA
           ,x"1001" -- 5DCC
           ,x"0559" -- 5DCE
           ,x"c809" -- 5DD0
           ,x"f076" -- 5DD2
           ,x"c820" -- 5DD4
           ,x"edd8" -- 5DD6
           ,x"f078" -- 5DD8
           ,x"0420" -- 5DDA
           ,x"137a" -- 5DDC
           ,x"0460" -- 5DDE
           ,x"8116" -- 5DE0
           ,x"c060" -- 5DE2
           ,x"ed0e" -- 5DE4
           ,x"c0c1" -- 5DE6
           ,x"0221" -- 5DE8
           ,x"fff6" -- 5DEA
           ,x"c801" -- 5DEC
           ,x"f076" -- 5DEE
           ,x"0420" -- 5DF0
           ,x"160e" -- 5DF2
           ,x"c083" -- 5DF4
           ,x"0222" -- 5DF6
           ,x"fff8" -- 5DF8
           ,x"a483" -- 5DFA
           ,x"c832" -- 5DFC
           ,x"edd2" -- 5DFE
           ,x"a483" -- 5E00
           ,x"c832" -- 5E02
           ,x"edd4" -- 5E04
           ,x"c820" -- 5E06
           ,x"f078" -- 5E08
           ,x"edd6" -- 5E0A
           ,x"6812" -- 5E0C
           ,x"edd6" -- 5E0E
           ,x"c820" -- 5E10
           ,x"f078" -- 5E12
           ,x"edd8" -- 5E14
           ,x"020e" -- 5E16
           ,x"aebe" -- 5E18
           ,x"020d" -- 5E1A
           ,x"efa8" -- 5E1C
           ,x"02cf" -- 5E1E
           ,x"0223" -- 5E20
           ,x"fff6" -- 5E22
           ,x"8813" -- 5E24
           ,x"c840" -- 5E26
           ,x"1302" -- 5E28
           ,x"0460" -- 5E2A
           ,x"8116" -- 5E2C
           ,x"0380" -- 5E2E
           ,x"0420" -- 5E30
           ,x"1744" -- 5E32
           ,x"0460" -- 5E34
           ,x"8116" -- 5E36
           ,x"4a00" -- 5E38
           ,x"c838" -- 5E3A
           ,x"4600" -- 5E3C
           ,x"c83c" -- 5E3E
           ,x"a5a5" -- 5E40
           ,x"457a" -- 5E42
           ,x"1200" -- 5E44
           ,x"0000" -- 5E46
           ,x"00f0" -- 5E48
           ,x"007f" -- 5E4A
           ,x"1331" -- 5E4C
           ,x"1b3c" -- 5E4E
           ,x"0d0a" -- 5E50
           ,x"2d2d" -- 5E52
           ,x"2054" -- 5E54
           ,x"4d53" -- 5E56
           ,x"2039" -- 5E58
           ,x"3939" -- 5E5A
           ,x"3520" -- 5E5C
           ,x"4272" -- 5E5E
           ,x"6561" -- 5E60
           ,x"6462" -- 5E62
           ,x"6f61" -- 5E64
           ,x"7264" -- 5E66
           ,x"2042" -- 5E68
           ,x"4153" -- 5E6A
           ,x"4943" -- 5E6C
           ,x"2052" -- 5E6E
           ,x"6576" -- 5E70
           ,x"2e20" -- 5E72
           ,x"312e" -- 5E74
           ,x"3120" -- 5E76
           ,x"2d2d" -- 5E78
           ,x"0d0a" -- 5E7A
           ,x"5b50" -- 5E7C
           ,x"6f72" -- 5E7E
           ,x"7465" -- 5E80
           ,x"6420" -- 5E82
           ,x"6672" -- 5E84
           ,x"6f6d" -- 5E86
           ,x"2043" -- 5E88
           ,x"6f72" -- 5E8A
           ,x"7465" -- 5E8C
           ,x"7820" -- 5E8E
           ,x"4241" -- 5E90
           ,x"5349" -- 5E92
           ,x"4320" -- 5E94
           ,x"2843" -- 5E96
           ,x"2931" -- 5E98
           ,x"3938" -- 5E9A
           ,x"3220" -- 5E9C
           ,x"6279" -- 5E9E
           ,x"2053" -- 5EA0
           ,x"7475" -- 5EA2
           ,x"6172" -- 5EA4
           ,x"7420" -- 5EA6
           ,x"436f" -- 5EA8
           ,x"6e6e" -- 5EAA
           ,x"6572" -- 5EAC
           ,x"5d0d" -- 5EAE
           ,x"0a0d" -- 5EB0
           ,x"0a2a" -- 5EB2
           ,x"5265" -- 5EB4
           ,x"6164" -- 5EB6
           ,x"790d" -- 5EB8
           ,x"0a00" -- 5EBA
           ,x"202a" -- 5EBC
           ,x"2ae0" -- 5EBE
           ,x"3f0d" -- 5EC0
           ,x"0a41" -- 5EC2
           ,x"7574" -- 5EC4
           ,x"6f2d" -- 5EC6
           ,x"5275" -- 5EC8
           ,x"6e20" -- 5ECA
           ,x"3f20" -- 5ECC
           ,x"2859" -- 5ECE
           ,x"2f4e" -- 5ED0
           ,x"29e0" -- 5ED2
           ,x"0d0a" -- 5ED4
           ,x"2a2a" -- 5ED6
           ,x"e03f" -- 5ED8
           ,x"3f20" -- 5EDA
           ,x"003a" -- 5EDC
           ,x"2000" -- 5EDE
           ,x"403e" -- 5EE0
           ,x"496e" -- 5EE2
           ,x"7661" -- 5EE4
           ,x"6c69" -- 5EE6
           ,x"6420" -- 5EE8
           ,x"6164" -- 5EEA
           ,x"6472" -- 5EEC
           ,x"6573" -- 5EEE
           ,x"8d00" -- 5EF0
           ,x"0000" -- 5EF2
           ,x"0000" -- 5EF4
           ,x"0000" -- 5EF6
           ,x"0000" -- 5EF8
           ,x"0000" -- 5EFA
           ,x"0000" -- 5EFC
           ,x"0000" -- 5EFE
           ,x"0000" -- 5F00
           ,x"0000" -- 5F02
           ,x"0000" -- 5F04
           ,x"0000" -- 5F06
           ,x"0000" -- 5F08
           ,x"0000" -- 5F0A
           ,x"0000" -- 5F0C
           ,x"0000" -- 5F0E
           ,x"0000" -- 5F10
           ,x"0000" -- 5F12
           ,x"0000" -- 5F14
           ,x"0000" -- 5F16
           ,x"0000" -- 5F18
           ,x"0000" -- 5F1A
           ,x"0000" -- 5F1C
           ,x"0000" -- 5F1E
           ,x"0000" -- 5F20
           ,x"0000" -- 5F22
           ,x"0000" -- 5F24
           ,x"0000" -- 5F26
           ,x"0000" -- 5F28
           ,x"0000" -- 5F2A
           ,x"0000" -- 5F2C
           ,x"0000" -- 5F2E
           ,x"0000" -- 5F30
           ,x"0000" -- 5F32
           ,x"0000" -- 5F34
           ,x"0000" -- 5F36
           ,x"0000" -- 5F38
           ,x"0000" -- 5F3A
           ,x"0000" -- 5F3C
           ,x"0000" -- 5F3E
           ,x"0000" -- 5F40
           ,x"0000" -- 5F42
           ,x"0000" -- 5F44
           ,x"0000" -- 5F46
           ,x"0000" -- 5F48
           ,x"0000" -- 5F4A
           ,x"0000" -- 5F4C
           ,x"0000" -- 5F4E
           ,x"0000" -- 5F50
           ,x"0000" -- 5F52
           ,x"0000" -- 5F54
           ,x"0000" -- 5F56
           ,x"0000" -- 5F58
           ,x"0000" -- 5F5A
           ,x"0000" -- 5F5C
           ,x"0000" -- 5F5E
           ,x"0000" -- 5F60
           ,x"0000" -- 5F62
           ,x"0000" -- 5F64
           ,x"0000" -- 5F66
           ,x"0000" -- 5F68
           ,x"0000" -- 5F6A
           ,x"0000" -- 5F6C
           ,x"0000" -- 5F6E
           ,x"0000" -- 5F70
           ,x"0000" -- 5F72
           ,x"0000" -- 5F74
           ,x"0000" -- 5F76
           ,x"0000" -- 5F78
           ,x"0000" -- 5F7A
           ,x"0000" -- 5F7C
           ,x"0000" -- 5F7E
           ,x"0000" -- 5F80
           ,x"0000" -- 5F82
           ,x"0000" -- 5F84
           ,x"0000" -- 5F86
           ,x"0000" -- 5F88
           ,x"0000" -- 5F8A
           ,x"0000" -- 5F8C
           ,x"0000" -- 5F8E
           ,x"0000" -- 5F90
           ,x"0000" -- 5F92
           ,x"0000" -- 5F94
           ,x"0000" -- 5F96
           ,x"0000" -- 5F98
           ,x"0000" -- 5F9A
           ,x"0000" -- 5F9C
           ,x"0000" -- 5F9E
           ,x"0000" -- 5FA0
           ,x"0000" -- 5FA2
           ,x"0000" -- 5FA4
           ,x"0000" -- 5FA6
           ,x"0000" -- 5FA8
           ,x"0000" -- 5FAA
           ,x"0000" -- 5FAC
           ,x"0000" -- 5FAE
           ,x"0000" -- 5FB0
           ,x"0000" -- 5FB2
           ,x"0000" -- 5FB4
           ,x"0000" -- 5FB6
           ,x"0000" -- 5FB8
           ,x"0000" -- 5FBA
           ,x"0000" -- 5FBC
           ,x"0000" -- 5FBE
           ,x"0000" -- 5FC0
           ,x"0000" -- 5FC2
           ,x"0000" -- 5FC4
           ,x"0000" -- 5FC6
           ,x"0000" -- 5FC8
           ,x"0000" -- 5FCA
           ,x"0000" -- 5FCC
           ,x"0000" -- 5FCE
           ,x"0000" -- 5FD0
           ,x"0000" -- 5FD2
           ,x"0000" -- 5FD4
           ,x"0000" -- 5FD6
           ,x"0000" -- 5FD8
           ,x"0000" -- 5FDA
           ,x"0000" -- 5FDC
           ,x"0000" -- 5FDE
           ,x"0000" -- 5FE0
           ,x"0000" -- 5FE2
           ,x"0000" -- 5FE4
           ,x"0000" -- 5FE6
           ,x"0000" -- 5FE8
           ,x"0000" -- 5FEA
           ,x"0000" -- 5FEC
           ,x"0000" -- 5FEE
           ,x"0000" -- 5FF0
           ,x"0000" -- 5FF2
           ,x"0000" -- 5FF4
           ,x"0000" -- 5FF6
           ,x"0000" -- 5FF8
           ,x"0000" -- 5FFA
           ,x"0000" -- 5FFC
           ,x"0000" -- 5FFE
           ,x"0000" -- 6000
           ,x"0000" -- 6002
           ,x"0000" -- 6004
           ,x"0000" -- 6006
           ,x"0000" -- 6008
           ,x"0000" -- 600A
           ,x"0000" -- 600C
           ,x"0000" -- 600E
           ,x"0000" -- 6010
           ,x"0000" -- 6012
           ,x"0000" -- 6014
           ,x"0000" -- 6016
           ,x"0000" -- 6018
           ,x"0000" -- 601A
           ,x"0000" -- 601C
           ,x"0000" -- 601E
           ,x"0000" -- 6020
           ,x"0000" -- 6022
           ,x"0000" -- 6024
           ,x"0000" -- 6026
           ,x"0000" -- 6028
           ,x"0000" -- 602A
           ,x"0000" -- 602C
           ,x"0000" -- 602E
           ,x"0000" -- 6030
           ,x"0000" -- 6032
           ,x"0000" -- 6034
           ,x"0000" -- 6036
           ,x"0000" -- 6038
           ,x"0000" -- 603A
           ,x"0000" -- 603C
           ,x"0000" -- 603E
           ,x"0000" -- 6040
           ,x"0000" -- 6042
           ,x"0000" -- 6044
           ,x"0000" -- 6046
           ,x"0000" -- 6048
           ,x"0000" -- 604A
           ,x"0000" -- 604C
           ,x"0000" -- 604E
           ,x"0000" -- 6050
           ,x"0000" -- 6052
           ,x"0000" -- 6054
           ,x"0000" -- 6056
           ,x"0000" -- 6058
           ,x"0000" -- 605A
           ,x"0000" -- 605C
           ,x"0000" -- 605E
           ,x"0000" -- 6060
           ,x"0000" -- 6062
           ,x"0000" -- 6064
           ,x"0000" -- 6066
           ,x"0000" -- 6068
           ,x"0000" -- 606A
           ,x"0000" -- 606C
           ,x"0000" -- 606E
           ,x"0000" -- 6070
           ,x"0000" -- 6072
           ,x"0000" -- 6074
           ,x"0000" -- 6076
           ,x"0000" -- 6078
           ,x"0000" -- 607A
           ,x"0000" -- 607C
           ,x"0000" -- 607E
           ,x"0000" -- 6080
           ,x"0000" -- 6082
           ,x"0000" -- 6084
           ,x"0000" -- 6086
           ,x"0000" -- 6088
           ,x"0000" -- 608A
           ,x"0000" -- 608C
           ,x"0000" -- 608E
           ,x"0000" -- 6090
           ,x"0000" -- 6092
           ,x"0000" -- 6094
           ,x"0000" -- 6096
           ,x"0000" -- 6098
           ,x"0000" -- 609A
           ,x"0000" -- 609C
           ,x"0000" -- 609E
           ,x"0000" -- 60A0
           ,x"0000" -- 60A2
           ,x"0000" -- 60A4
           ,x"0000" -- 60A6
           ,x"0000" -- 60A8
           ,x"0000" -- 60AA
           ,x"0000" -- 60AC
           ,x"0000" -- 60AE
           ,x"0000" -- 60B0
           ,x"0000" -- 60B2
           ,x"0000" -- 60B4
           ,x"0000" -- 60B6
           ,x"0000" -- 60B8
           ,x"0000" -- 60BA
           ,x"0000" -- 60BC
           ,x"0000" -- 60BE
           ,x"0000" -- 60C0
           ,x"0000" -- 60C2
           ,x"0000" -- 60C4
           ,x"0000" -- 60C6
           ,x"0000" -- 60C8
           ,x"0000" -- 60CA
           ,x"0000" -- 60CC
           ,x"0000" -- 60CE
           ,x"0000" -- 60D0
           ,x"0000" -- 60D2
           ,x"0000" -- 60D4
           ,x"0000" -- 60D6
           ,x"0000" -- 60D8
           ,x"0000" -- 60DA
           ,x"0000" -- 60DC
           ,x"0000" -- 60DE
           ,x"0000" -- 60E0
           ,x"0000" -- 60E2
           ,x"0000" -- 60E4
           ,x"0000" -- 60E6
           ,x"0000" -- 60E8
           ,x"0000" -- 60EA
           ,x"0000" -- 60EC
           ,x"0000" -- 60EE
           ,x"0000" -- 60F0
           ,x"0000" -- 60F2
           ,x"0000" -- 60F4
           ,x"0000" -- 60F6
           ,x"0000" -- 60F8
           ,x"0000" -- 60FA
           ,x"0000" -- 60FC
           ,x"0000" -- 60FE
           ,x"0000" -- 6100
           ,x"0000" -- 6102
           ,x"0000" -- 6104
           ,x"0000" -- 6106
           ,x"0000" -- 6108
           ,x"0000" -- 610A
           ,x"0000" -- 610C
           ,x"0000" -- 610E
           ,x"0000" -- 6110
           ,x"0000" -- 6112
           ,x"0000" -- 6114
           ,x"0000" -- 6116
           ,x"0000" -- 6118
           ,x"0000" -- 611A
           ,x"0000" -- 611C
           ,x"0000" -- 611E
           ,x"0000" -- 6120
           ,x"0000" -- 6122
           ,x"0000" -- 6124
           ,x"0000" -- 6126
           ,x"0000" -- 6128
           ,x"0000" -- 612A
           ,x"0000" -- 612C
           ,x"0000" -- 612E
           ,x"0000" -- 6130
           ,x"0000" -- 6132
           ,x"0000" -- 6134
           ,x"0000" -- 6136
           ,x"0000" -- 6138
           ,x"0000" -- 613A
           ,x"0000" -- 613C
           ,x"0000" -- 613E
           ,x"0000" -- 6140
           ,x"0000" -- 6142
           ,x"0000" -- 6144
           ,x"0000" -- 6146
           ,x"0000" -- 6148
           ,x"0000" -- 614A
           ,x"0000" -- 614C
           ,x"0000" -- 614E
           ,x"0000" -- 6150
           ,x"0000" -- 6152
           ,x"0000" -- 6154
           ,x"0000" -- 6156
           ,x"0000" -- 6158
           ,x"0000" -- 615A
           ,x"0000" -- 615C
           ,x"0000" -- 615E
           ,x"0000" -- 6160
           ,x"0000" -- 6162
           ,x"0000" -- 6164
           ,x"0000" -- 6166
           ,x"0000" -- 6168
           ,x"0000" -- 616A
           ,x"0000" -- 616C
           ,x"0000" -- 616E
           ,x"0000" -- 6170
           ,x"0000" -- 6172
           ,x"0000" -- 6174
           ,x"0000" -- 6176
           ,x"0000" -- 6178
           ,x"0000" -- 617A
           ,x"0000" -- 617C
           ,x"0000" -- 617E
           ,x"0000" -- 6180
           ,x"0000" -- 6182
           ,x"0000" -- 6184
           ,x"0000" -- 6186
           ,x"0000" -- 6188
           ,x"0000" -- 618A
           ,x"0000" -- 618C
           ,x"0000" -- 618E
           ,x"0000" -- 6190
           ,x"0000" -- 6192
           ,x"0000" -- 6194
           ,x"0000" -- 6196
           ,x"0000" -- 6198
           ,x"0000" -- 619A
           ,x"0000" -- 619C
           ,x"0000" -- 619E
           ,x"0000" -- 61A0
           ,x"0000" -- 61A2
           ,x"0000" -- 61A4
           ,x"0000" -- 61A6
           ,x"0000" -- 61A8
           ,x"0000" -- 61AA
           ,x"0000" -- 61AC
           ,x"0000" -- 61AE
           ,x"0000" -- 61B0
           ,x"0000" -- 61B2
           ,x"0000" -- 61B4
           ,x"0000" -- 61B6
           ,x"0000" -- 61B8
           ,x"0000" -- 61BA
           ,x"0000" -- 61BC
           ,x"0000" -- 61BE
           ,x"0000" -- 61C0
           ,x"0000" -- 61C2
           ,x"0000" -- 61C4
           ,x"0000" -- 61C6
           ,x"0000" -- 61C8
           ,x"0000" -- 61CA
           ,x"0000" -- 61CC
           ,x"0000" -- 61CE
           ,x"0000" -- 61D0
           ,x"0000" -- 61D2
           ,x"0000" -- 61D4
           ,x"0000" -- 61D6
           ,x"0000" -- 61D8
           ,x"0000" -- 61DA
           ,x"0000" -- 61DC
           ,x"0000" -- 61DE
           ,x"0000" -- 61E0
           ,x"0000" -- 61E2
           ,x"0000" -- 61E4
           ,x"0000" -- 61E6
           ,x"0000" -- 61E8
           ,x"0000" -- 61EA
           ,x"0000" -- 61EC
           ,x"0000" -- 61EE
           ,x"0000" -- 61F0
           ,x"0000" -- 61F2
           ,x"0000" -- 61F4
           ,x"0000" -- 61F6
           ,x"0000" -- 61F8
           ,x"0000" -- 61FA
           ,x"0000" -- 61FC
           ,x"0000" -- 61FE
           ,x"0000" -- 6200
           ,x"0000" -- 6202
           ,x"0000" -- 6204
           ,x"0000" -- 6206
           ,x"0000" -- 6208
           ,x"0000" -- 620A
           ,x"0000" -- 620C
           ,x"0000" -- 620E
           ,x"0000" -- 6210
           ,x"0000" -- 6212
           ,x"0000" -- 6214
           ,x"0000" -- 6216
           ,x"0000" -- 6218
           ,x"0000" -- 621A
           ,x"0000" -- 621C
           ,x"0000" -- 621E
           ,x"0000" -- 6220
           ,x"0000" -- 6222
           ,x"0000" -- 6224
           ,x"0000" -- 6226
           ,x"0000" -- 6228
           ,x"0000" -- 622A
           ,x"0000" -- 622C
           ,x"0000" -- 622E
           ,x"0000" -- 6230
           ,x"0000" -- 6232
           ,x"0000" -- 6234
           ,x"0000" -- 6236
           ,x"0000" -- 6238
           ,x"0000" -- 623A
           ,x"0000" -- 623C
           ,x"0000" -- 623E
           ,x"0000" -- 6240
           ,x"0000" -- 6242
           ,x"0000" -- 6244
           ,x"0000" -- 6246
           ,x"0000" -- 6248
           ,x"0000" -- 624A
           ,x"0000" -- 624C
           ,x"0000" -- 624E
           ,x"0000" -- 6250
           ,x"0000" -- 6252
           ,x"0000" -- 6254
           ,x"0000" -- 6256
           ,x"0000" -- 6258
           ,x"0000" -- 625A
           ,x"0000" -- 625C
           ,x"0000" -- 625E
           ,x"0000" -- 6260
           ,x"0000" -- 6262
           ,x"0000" -- 6264
           ,x"0000" -- 6266
           ,x"0000" -- 6268
           ,x"0000" -- 626A
           ,x"0000" -- 626C
           ,x"0000" -- 626E
           ,x"0000" -- 6270
           ,x"0000" -- 6272
           ,x"0000" -- 6274
           ,x"0000" -- 6276
           ,x"0000" -- 6278
           ,x"0000" -- 627A
           ,x"0000" -- 627C
           ,x"0000" -- 627E
           ,x"0000" -- 6280
           ,x"0000" -- 6282
           ,x"0000" -- 6284
           ,x"0000" -- 6286
           ,x"0000" -- 6288
           ,x"eb0e" -- 628A
           ,x"ecfe" -- 628C
           ,x"ec4a" -- 628E
           ,x"ebfa" -- 6290
           ,x"eb8e" -- 6292
           ,x"02e0" -- 6294
           ,x"efa8" -- 6296
           ,x"0202" -- 6298
           ,x"efa8" -- 629A
           ,x"0642" -- 629C
           ,x"04d2" -- 629E
           ,x"0282" -- 62A0
           ,x"dab0" -- 62A2
           ,x"1bfb" -- 62A4
           ,x"0201" -- 62A6
           ,x"ed04" -- 62A8
           ,x"0205" -- 62AA
           ,x"cc8a" -- 62AC
           ,x"0222" -- 62AE
           ,x"000a" -- 62B0
           ,x"c802" -- 62B2
           ,x"8048" -- 62B4
           ,x"0202" -- 62B6
           ,x"deba" -- 62B8
           ,x"cc75" -- 62BA
           ,x"cc75" -- 62BC
           ,x"cc75" -- 62BE
           ,x"cc75" -- 62C0
           ,x"cc55" -- 62C2
           ,x"cc42" -- 62C4
           ,x"cc42" -- 62C6
           ,x"0201" -- 62C8
           ,x"d6ba" -- 62CA
           ,x"0202" -- 62CC
           ,x"d0ba" -- 62CE
           ,x"ccb1" -- 62D0
           ,x"0282" -- 62D2
           ,x"d4b0" -- 62D4
           ,x"1afc" -- 62D6
           ,x"020b" -- 62D8
           ,x"80ee" -- 62DA
           ,x"0460" -- 62DC
           ,x"8094" -- 62DE
           ,x"5359" -- 62E0
           ,x"5354" -- 62E2
           ,x"454d" -- 62E4
           ,x"2045" -- 62E6
           ,x"5252" -- 62E8
           ,x"4fae" -- 62EA
           ,x"5379" -- 62EC
           ,x"6e74" -- 62EE
           ,x"6178" -- 62F0
           ,x"2065" -- 62F2
           ,x"7272" -- 62F4
           ,x"6f8e" -- 62F6
           ,x"556e" -- 62F8
           ,x"6d61" -- 62FA
           ,x"7463" -- 62FC
           ,x"6865" -- 62FE
           ,x"6420" -- 6300
           ,x"6465" -- 6302
           ,x"6c69" -- 6304
           ,x"6d69" -- 6306
           ,x"7465" -- 6308
           ,x"8e49" -- 630A
           ,x"6e76" -- 630C
           ,x"616c" -- 630E
           ,x"6964" -- 6310
           ,x"206c" -- 6312
           ,x"696e" -- 6314
           ,x"6520" -- 6316
           ,x"6e75" -- 6318
           ,x"6d62" -- 631A
           ,x"658e" -- 631C
           ,x"496c" -- 631E
           ,x"6c65" -- 6320
           ,x"6761" -- 6322
           ,x"6c20" -- 6324
           ,x"7661" -- 6326
           ,x"7269" -- 6328
           ,x"6162" -- 632A
           ,x"6c65" -- 632C
           ,x"206e" -- 632E
           ,x"616d" -- 6330
           ,x"9b54" -- 6332
           ,x"6f6f" -- 6334
           ,x"206d" -- 6336
           ,x"616e" -- 6338
           ,x"7920" -- 633A
           ,x"7661" -- 633C
           ,x"7269" -- 633E
           ,x"6162" -- 6340
           ,x"6c65" -- 6342
           ,x"8d49" -- 6344
           ,x"6c6c" -- 6346
           ,x"6567" -- 6348
           ,x"616c" -- 634A
           ,x"2063" -- 634C
           ,x"6861" -- 634E
           ,x"7261" -- 6350
           ,x"6374" -- 6352
           ,x"658e" -- 6354
           ,x"4578" -- 6356
           ,x"7065" -- 6358
           ,x"6374" -- 635A
           ,x"696e" -- 635C
           ,x"6720" -- 635E
           ,x"6f70" -- 6360
           ,x"6572" -- 6362
           ,x"6174" -- 6364
           ,x"6f8e" -- 6366
           ,x"496c" -- 6368
           ,x"6c65" -- 636A
           ,x"6761" -- 636C
           ,x"6c20" -- 636E
           ,x"6675" -- 6370
           ,x"6e63" -- 6372
           ,x"7469" -- 6374
           ,x"6f6e" -- 6376
           ,x"206e" -- 6378
           ,x"616d" -- 637A
           ,x"9b49" -- 637C
           ,x"6c6c" -- 637E
           ,x"6567" -- 6380
           ,x"616c" -- 6382
           ,x"2066" -- 6384
           ,x"756e" -- 6386
           ,x"6374" -- 6388
           ,x"696f" -- 638A
           ,x"6e20" -- 638C
           ,x"6172" -- 638E
           ,x"6775" -- 6390
           ,x"6d65" -- 6392
           ,x"6e8c" -- 6394
           ,x"4f75" -- 6396
           ,x"7420" -- 6398
           ,x"6f66" -- 639A
           ,x"206d" -- 639C
           ,x"656d" -- 639E
           ,x"6f72" -- 63A0
           ,x"8753" -- 63A2
           ,x"7461" -- 63A4
           ,x"636b" -- 63A6
           ,x"206f" -- 63A8
           ,x"7665" -- 63AA
           ,x"7266" -- 63AC
           ,x"6c6f" -- 63AE
           ,x"8953" -- 63B0
           ,x"7461" -- 63B2
           ,x"636b" -- 63B4
           ,x"2075" -- 63B6
           ,x"6e64" -- 63B8
           ,x"6572" -- 63BA
           ,x"666c" -- 63BC
           ,x"6f89" -- 63BE
           ,x"4e6f" -- 63C0
           ,x"2073" -- 63C2
           ,x"7563" -- 63C4
           ,x"6820" -- 63C6
           ,x"6c69" -- 63C8
           ,x"6e65" -- 63CA
           ,x"206e" -- 63CC
           ,x"756d" -- 63CE
           ,x"6265" -- 63D0
           ,x"8e45" -- 63D2
           ,x"7870" -- 63D4
           ,x"6563" -- 63D6
           ,x"7469" -- 63D8
           ,x"6e67" -- 63DA
           ,x"2073" -- 63DC
           ,x"7472" -- 63DE
           ,x"696e" -- 63E0
           ,x"6720" -- 63E2
           ,x"7661" -- 63E4
           ,x"7269" -- 63E6
           ,x"6162" -- 63E8
           ,x"6c9b" -- 63EA
           ,x"496e" -- 63EC
           ,x"7661" -- 63EE
           ,x"6c69" -- 63F0
           ,x"6420" -- 63F2
           ,x"7363" -- 63F4
           ,x"7265" -- 63F6
           ,x"656e" -- 63F8
           ,x"2063" -- 63FA
           ,x"6f6d" -- 63FC
           ,x"6d61" -- 63FE
           ,x"6e9c" -- 6400
           ,x"4578" -- 6402
           ,x"7065" -- 6404
           ,x"6374" -- 6406
           ,x"696e" -- 6408
           ,x"6720" -- 640A
           ,x"6469" -- 640C
           ,x"6d65" -- 640E
           ,x"6e73" -- 6410
           ,x"696f" -- 6412
           ,x"6e65" -- 6414
           ,x"6420" -- 6416
           ,x"7661" -- 6418
           ,x"7269" -- 641A
           ,x"6162" -- 641C
           ,x"6c9b" -- 641E
           ,x"5375" -- 6420
           ,x"6273" -- 6422
           ,x"6372" -- 6424
           ,x"6970" -- 6426
           ,x"7420" -- 6428
           ,x"6f75" -- 642A
           ,x"7420" -- 642C
           ,x"6f66" -- 642E
           ,x"2072" -- 6430
           ,x"616e" -- 6432
           ,x"679b" -- 6434
           ,x"546f" -- 6436
           ,x"6f20" -- 6438
           ,x"6665" -- 643A
           ,x"7720" -- 643C
           ,x"7375" -- 643E
           ,x"6273" -- 6440
           ,x"6372" -- 6442
           ,x"6970" -- 6444
           ,x"748d" -- 6446
           ,x"546f" -- 6448
           ,x"6f20" -- 644A
           ,x"6d61" -- 644C
           ,x"6e79" -- 644E
           ,x"2073" -- 6450
           ,x"7562" -- 6452
           ,x"7363" -- 6454
           ,x"7269" -- 6456
           ,x"7074" -- 6458
           ,x"8d45" -- 645A
           ,x"7870" -- 645C
           ,x"6563" -- 645E
           ,x"7469" -- 6460
           ,x"6e67" -- 6462
           ,x"2073" -- 6464
           ,x"696d" -- 6466
           ,x"706c" -- 6468
           ,x"6520" -- 646A
           ,x"7661" -- 646C
           ,x"7269" -- 646E
           ,x"6162" -- 6470
           ,x"6c9b" -- 6472
           ,x"4578" -- 6474
           ,x"7065" -- 6476
           ,x"6374" -- 6478
           ,x"696e" -- 647A
           ,x"6720" -- 647C
           ,x"7661" -- 647E
           ,x"7269" -- 6480
           ,x"6162" -- 6482
           ,x"6c9b" -- 6484
           ,x"5265" -- 6486
           ,x"6164" -- 6488
           ,x"206f" -- 648A
           ,x"7574" -- 648C
           ,x"206f" -- 648E
           ,x"6620" -- 6490
           ,x"4461" -- 6492
           ,x"749f" -- 6494
           ,x"5265" -- 6496
           ,x"6164" -- 6498
           ,x"2026" -- 649A
           ,x"2044" -- 649C
           ,x"6174" -- 649E
           ,x"6120" -- 64A0
           ,x"7479" -- 64A2
           ,x"7065" -- 64A4
           ,x"7320" -- 64A6
           ,x"6469" -- 64A8
           ,x"6666" -- 64AA
           ,x"658e" -- 64AC
           ,x"5371" -- 64AE
           ,x"7561" -- 64B0
           ,x"7265" -- 64B2
           ,x"2072" -- 64B4
           ,x"6f6f" -- 64B6
           ,x"7420" -- 64B8
           ,x"6f66" -- 64BA
           ,x"206e" -- 64BC
           ,x"6567" -- 64BE
           ,x"6174" -- 64C0
           ,x"6976" -- 64C2
           ,x"6520" -- 64C4
           ,x"6e75" -- 64C6
           ,x"6d62" -- 64C8
           ,x"658e" -- 64CA
           ,x"4c6f" -- 64CC
           ,x"6720" -- 64CE
           ,x"6f66" -- 64D0
           ,x"206e" -- 64D2
           ,x"6f6e" -- 64D4
           ,x"2d70" -- 64D6
           ,x"6f73" -- 64D8
           ,x"6974" -- 64DA
           ,x"6976" -- 64DC
           ,x"6520" -- 64DE
           ,x"6e75" -- 64E0
           ,x"6d62" -- 64E2
           ,x"658e" -- 64E4
           ,x"4578" -- 64E6
           ,x"7072" -- 64E8
           ,x"6573" -- 64EA
           ,x"7369" -- 64EC
           ,x"6f6e" -- 64EE
           ,x"2074" -- 64F0
           ,x"6f6f" -- 64F2
           ,x"2063" -- 64F4
           ,x"6f6d" -- 64F6
           ,x"706c" -- 64F8
           ,x"6588" -- 64FA
           ,x"4469" -- 64FC
           ,x"7669" -- 64FE
           ,x"7369" -- 6500
           ,x"6f6e" -- 6502
           ,x"2062" -- 6504
           ,x"7920" -- 6506
           ,x"7a65" -- 6508
           ,x"7291" -- 650A
           ,x"466c" -- 650C
           ,x"6f61" -- 650E
           ,x"7469" -- 6510
           ,x"6e67" -- 6512
           ,x"2070" -- 6514
           ,x"6f69" -- 6516
           ,x"6e74" -- 6518
           ,x"206f" -- 651A
           ,x"7665" -- 651C
           ,x"7266" -- 651E
           ,x"6c6f" -- 6520
           ,x"8952" -- 6522
           ,x"616e" -- 6524
           ,x"6765" -- 6526
           ,x"2065" -- 6528
           ,x"7272" -- 652A
           ,x"6f8e" -- 652C
           ,x"4d69" -- 652E
           ,x"7373" -- 6530
           ,x"696e" -- 6532
           ,x"6720" -- 6534
           ,x"4e45" -- 6536
           ,x"58ac" -- 6538
           ,x"4d69" -- 653A
           ,x"7373" -- 653C
           ,x"696e" -- 653E
           ,x"6720" -- 6540
           ,x"464f" -- 6542
           ,x"ae45" -- 6544
           ,x"5850" -- 6546
           ,x"2068" -- 6548
           ,x"6173" -- 654A
           ,x"2069" -- 654C
           ,x"6e76" -- 654E
           ,x"616c" -- 6550
           ,x"6964" -- 6552
           ,x"2061" -- 6554
           ,x"7267" -- 6556
           ,x"756d" -- 6558
           ,x"656e" -- 655A
           ,x"8c55" -- 655C
           ,x"6e6e" -- 655E
           ,x"6f72" -- 6560
           ,x"6d61" -- 6562
           ,x"6c69" -- 6564
           ,x"7365" -- 6566
           ,x"6420" -- 6568
           ,x"6e75" -- 656A
           ,x"6d62" -- 656C
           ,x"658e" -- 656E
           ,x"5061" -- 6570
           ,x"7261" -- 6572
           ,x"6d65" -- 6574
           ,x"7465" -- 6576
           ,x"7220" -- 6578
           ,x"6572" -- 657A
           ,x"726f" -- 657C
           ,x"8e4d" -- 657E
           ,x"6973" -- 6580
           ,x"7369" -- 6582
           ,x"6e67" -- 6584
           ,x"2061" -- 6586
           ,x"7373" -- 6588
           ,x"6967" -- 658A
           ,x"6e6d" -- 658C
           ,x"656e" -- 658E
           ,x"7420" -- 6590
           ,x"6f70" -- 6592
           ,x"6572" -- 6594
           ,x"6174" -- 6596
           ,x"6f8e" -- 6598
           ,x"496c" -- 659A
           ,x"6c65" -- 659C
           ,x"6761" -- 659E
           ,x"6c20" -- 65A0
           ,x"6465" -- 65A2
           ,x"6c69" -- 65A4
           ,x"6d69" -- 65A6
           ,x"7465" -- 65A8
           ,x"8e55" -- 65AA
           ,x"6e64" -- 65AC
           ,x"6566" -- 65AE
           ,x"696e" -- 65B0
           ,x"6564" -- 65B2
           ,x"2066" -- 65B4
           ,x"756e" -- 65B6
           ,x"6374" -- 65B8
           ,x"696f" -- 65BA
           ,x"9255" -- 65BC
           ,x"6e64" -- 65BE
           ,x"696d" -- 65C0
           ,x"656e" -- 65C2
           ,x"7369" -- 65C4
           ,x"6f6e" -- 65C6
           ,x"6564" -- 65C8
           ,x"2076" -- 65CA
           ,x"6172" -- 65CC
           ,x"6961" -- 65CE
           ,x"626c" -- 65D0
           ,x"9b55" -- 65D2
           ,x"6e64" -- 65D4
           ,x"6566" -- 65D6
           ,x"696e" -- 65D8
           ,x"6564" -- 65DA
           ,x"2076" -- 65DC
           ,x"6172" -- 65DE
           ,x"6961" -- 65E0
           ,x"626c" -- 65E2
           ,x"9b45" -- 65E4
           ,x"7874" -- 65E6
           ,x"6572" -- 65E8
           ,x"6e61" -- 65EA
           ,x"6c20" -- 65EC
           ,x"636f" -- 65EE
           ,x"6d6d" -- 65F0
           ,x"616e" -- 65F2
           ,x"6420" -- 65F4
           ,x"6e6f" -- 65F6
           ,x"7420" -- 65F8
           ,x"666f" -- 65FA
           ,x"756e" -- 65FC
           ,x"9c49" -- 65FE
           ,x"6e76" -- 6600
           ,x"616c" -- 6602
           ,x"6964" -- 6604
           ,x"2064" -- 6606
           ,x"6576" -- 6608
           ,x"6963" -- 660A
           ,x"6520" -- 660C
           ,x"6e75" -- 660E
           ,x"6d62" -- 6610
           ,x"658e" -- 6612
           ,x"496c" -- 6614
           ,x"6c65" -- 6616
           ,x"6761" -- 6618
           ,x"6c20" -- 661A
           ,x"696e" -- 661C
           ,x"2063" -- 661E
           ,x"7572" -- 6620
           ,x"7265" -- 6622
           ,x"6e74" -- 6624
           ,x"206d" -- 6626
           ,x"6f64" -- 6628
           ,x"9b43" -- 662A
           ,x"6f6d" -- 662C
           ,x"6d61" -- 662E
           ,x"6e64" -- 6630
           ,x"206e" -- 6632
           ,x"6f74" -- 6634
           ,x"2073" -- 6636
           ,x"7570" -- 6638
           ,x"706f" -- 663A
           ,x"7274" -- 663C
           ,x"659c" -- 663E
           ,x"492f" -- 6640
           ,x"4f20" -- 6642
           ,x"6572" -- 6644
           ,x"726f" -- 6646
           ,x"7220" -- 6648
           ,x"636f" -- 664A
           ,x"6465" -- 664C
           ,x"2000" -- 664E
           ,x"ef00" -- 6650
           ,x"d054" -- 6652
           ,x"8289" -- 6654
           ,x"1b06" -- 6656
           ,x"d039" -- 6658
           ,x"9800" -- 665A
           ,x"c0e4" -- 665C
           ,x"1a03" -- 665E
           ,x"2f00" -- 6660
           ,x"10f8" -- 6662
           ,x"0380" -- 6664
           ,x"06a0" -- 6666
           ,x"872c" -- 6668
           ,x"0909" -- 666A
           ,x"0e08" -- 666C
           ,x"130a" -- 666E
           ,x"150b" -- 6670
           ,x"1a0c" -- 6672
           ,x"240d" -- 6674
           ,x"1d1e" -- 6676
           ,x"0000" -- 6678
           ,x"10ec" -- 667A
           ,x"2fa0" -- 667C
           ,x"d082" -- 667E
           ,x"10e9" -- 6680
           ,x"1b5b" -- 6682
           ,x"4300" -- 6684
           ,x"2fa0" -- 6686
           ,x"d08c" -- 6688
           ,x"10e4" -- 668A
           ,x"1b5b" -- 668C
           ,x"4400" -- 668E
           ,x"2f00" -- 6690
           ,x"10e0" -- 6692
           ,x"2fa0" -- 6694
           ,x"d09a" -- 6696
           ,x"10dd" -- 6698
           ,x"1b5b" -- 669A
           ,x"4100" -- 669C
           ,x"2fa0" -- 669E
           ,x"d0aa" -- 66A0
           ,x"10d8" -- 66A2
           ,x"2fa0" -- 66A4
           ,x"d0ae" -- 66A6
           ,x"10d5" -- 66A8
           ,x"1b5b" -- 66AA
           ,x"324a" -- 66AC
           ,x"1b5b" -- 66AE
           ,x"4800" -- 66B0
           ,x"2f00" -- 66B2
           ,x"04e0" -- 66B4
           ,x"ed34" -- 66B6
           ,x"10cd" -- 66B8
           ,x"0000" -- 66BA
           ,x"0000" -- 66BC
           ,x"0000" -- 66BE
           ,x"0000" -- 66C0
           ,x"0000" -- 66C2
           ,x"0000" -- 66C4
           ,x"0000" -- 66C6
           ,x"0000" -- 66C8
           ,x"0000" -- 66CA
           ,x"0000" -- 66CC
           ,x"0000" -- 66CE
           ,x"0000" -- 66D0
           ,x"0000" -- 66D2
           ,x"0000" -- 66D4
           ,x"0000" -- 66D6
           ,x"0000" -- 66D8
           ,x"0000" -- 66DA
           ,x"0000" -- 66DC
           ,x"0000" -- 66DE
           ,x"0000" -- 66E0
           ,x"0000" -- 66E2
           ,x"0000" -- 66E4
           ,x"0000" -- 66E6
           ,x"0000" -- 66E8
           ,x"0000" -- 66EA
           ,x"0000" -- 66EC
           ,x"0000" -- 66EE
           ,x"0000" -- 66F0
           ,x"0000" -- 66F2
           ,x"0000" -- 66F4
           ,x"0000" -- 66F6
           ,x"0000" -- 66F8
           ,x"0000" -- 66FA
           ,x"0000" -- 66FC
           ,x"0000" -- 66FE
           ,x"0000" -- 6700
           ,x"0000" -- 6702
           ,x"0000" -- 6704
           ,x"0000" -- 6706
           ,x"0000" -- 6708
           ,x"0000" -- 670A
           ,x"0000" -- 670C
           ,x"0000" -- 670E
           ,x"0000" -- 6710
           ,x"0000" -- 6712
           ,x"0000" -- 6714
           ,x"0000" -- 6716
           ,x"0000" -- 6718
           ,x"0000" -- 671A
           ,x"0000" -- 671C
           ,x"0000" -- 671E
           ,x"0000" -- 6720
           ,x"0000" -- 6722
           ,x"0000" -- 6724
           ,x"0000" -- 6726
           ,x"0000" -- 6728
           ,x"0000" -- 672A
           ,x"0000" -- 672C
           ,x"0000" -- 672E
           ,x"0000" -- 6730
           ,x"0000" -- 6732
           ,x"0000" -- 6734
           ,x"0000" -- 6736
           ,x"0000" -- 6738
           ,x"0000" -- 673A
           ,x"0000" -- 673C
           ,x"0000" -- 673E
           ,x"0000" -- 6740
           ,x"0000" -- 6742
           ,x"0000" -- 6744
           ,x"0000" -- 6746
           ,x"0000" -- 6748
           ,x"0000" -- 674A
           ,x"0000" -- 674C
           ,x"0000" -- 674E
           ,x"0000" -- 6750
           ,x"0000" -- 6752
           ,x"0000" -- 6754
           ,x"0000" -- 6756
           ,x"0000" -- 6758
           ,x"0000" -- 675A
           ,x"0000" -- 675C
           ,x"0000" -- 675E
           ,x"0000" -- 6760
           ,x"0000" -- 6762
           ,x"0000" -- 6764
           ,x"0000" -- 6766
           ,x"0000" -- 6768
           ,x"0000" -- 676A
           ,x"0000" -- 676C
           ,x"0000" -- 676E
           ,x"0000" -- 6770
           ,x"0000" -- 6772
           ,x"0000" -- 6774
           ,x"0000" -- 6776
           ,x"0000" -- 6778
           ,x"0000" -- 677A
           ,x"0000" -- 677C
           ,x"0000" -- 677E
           ,x"0000" -- 6780
           ,x"0000" -- 6782
           ,x"0000" -- 6784
           ,x"0000" -- 6786
           ,x"0000" -- 6788
           ,x"0000" -- 678A
           ,x"0000" -- 678C
           ,x"0000" -- 678E
           ,x"0000" -- 6790
           ,x"0000" -- 6792
           ,x"0000" -- 6794
           ,x"0000" -- 6796
           ,x"0000" -- 6798
           ,x"0000" -- 679A
           ,x"0000" -- 679C
           ,x"0000" -- 679E
           ,x"0000" -- 67A0
           ,x"0000" -- 67A2
           ,x"0000" -- 67A4
           ,x"0000" -- 67A6
           ,x"0000" -- 67A8
           ,x"0000" -- 67AA
           ,x"0000" -- 67AC
           ,x"0000" -- 67AE
           ,x"0000" -- 67B0
           ,x"0000" -- 67B2
           ,x"0000" -- 67B4
           ,x"0000" -- 67B6
           ,x"0000" -- 67B8
           ,x"0000" -- 67BA
           ,x"0000" -- 67BC
           ,x"0000" -- 67BE
           ,x"0000" -- 67C0
           ,x"0000" -- 67C2
           ,x"0000" -- 67C4
           ,x"0000" -- 67C6
           ,x"0000" -- 67C8
           ,x"0000" -- 67CA
           ,x"0000" -- 67CC
           ,x"0000" -- 67CE
           ,x"0000" -- 67D0
           ,x"0000" -- 67D2
           ,x"0000" -- 67D4
           ,x"0000" -- 67D6
           ,x"0000" -- 67D8
           ,x"0000" -- 67DA
           ,x"0000" -- 67DC
           ,x"0000" -- 67DE
           ,x"0000" -- 67E0
           ,x"0000" -- 67E2
           ,x"0000" -- 67E4
           ,x"0000" -- 67E6
           ,x"0000" -- 67E8
           ,x"0000" -- 67EA
           ,x"0000" -- 67EC
           ,x"0000" -- 67EE
           ,x"0000" -- 67F0
           ,x"0000" -- 67F2
           ,x"0000" -- 67F4
           ,x"0000" -- 67F6
           ,x"0000" -- 67F8
           ,x"0000" -- 67FA
           ,x"0000" -- 67FC
           ,x"0000" -- 67FE
           ,x"0000" -- 6800
           ,x"0000" -- 6802
           ,x"0000" -- 6804
           ,x"0000" -- 6806
           ,x"0000" -- 6808
           ,x"0000" -- 680A
           ,x"0000" -- 680C
           ,x"0000" -- 680E
           ,x"0000" -- 6810
           ,x"0000" -- 6812
           ,x"0000" -- 6814
           ,x"0000" -- 6816
           ,x"0000" -- 6818
           ,x"0000" -- 681A
           ,x"0000" -- 681C
           ,x"0000" -- 681E
           ,x"0000" -- 6820
           ,x"0000" -- 6822
           ,x"0000" -- 6824
           ,x"0000" -- 6826
           ,x"0000" -- 6828
           ,x"0000" -- 682A
           ,x"0000" -- 682C
           ,x"0000" -- 682E
           ,x"0000" -- 6830
           ,x"0000" -- 6832
           ,x"0000" -- 6834
           ,x"0000" -- 6836
           ,x"0000" -- 6838
           ,x"0000" -- 683A
           ,x"0000" -- 683C
           ,x"0000" -- 683E
           ,x"0000" -- 6840
           ,x"0000" -- 6842
           ,x"0000" -- 6844
           ,x"0000" -- 6846
           ,x"0000" -- 6848
           ,x"0000" -- 684A
           ,x"0000" -- 684C
           ,x"0000" -- 684E
           ,x"0000" -- 6850
           ,x"0000" -- 6852
           ,x"0000" -- 6854
           ,x"0000" -- 6856
           ,x"0000" -- 6858
           ,x"0000" -- 685A
           ,x"0000" -- 685C
           ,x"0000" -- 685E
           ,x"0000" -- 6860
           ,x"0000" -- 6862
           ,x"0000" -- 6864
           ,x"0000" -- 6866
           ,x"0000" -- 6868
           ,x"0000" -- 686A
           ,x"0000" -- 686C
           ,x"0000" -- 686E
           ,x"0000" -- 6870
           ,x"0000" -- 6872
           ,x"0000" -- 6874
           ,x"0000" -- 6876
           ,x"0000" -- 6878
           ,x"0000" -- 687A
           ,x"0000" -- 687C
           ,x"0000" -- 687E
           ,x"0000" -- 6880
           ,x"0000" -- 6882
           ,x"0000" -- 6884
           ,x"0000" -- 6886
           ,x"0000" -- 6888
           ,x"0000" -- 688A
           ,x"0000" -- 688C
           ,x"0000" -- 688E
           ,x"0000" -- 6890
           ,x"0000" -- 6892
           ,x"0000" -- 6894
           ,x"0000" -- 6896
           ,x"0000" -- 6898
           ,x"0000" -- 689A
           ,x"0000" -- 689C
           ,x"0000" -- 689E
           ,x"0000" -- 68A0
           ,x"0000" -- 68A2
           ,x"0000" -- 68A4
           ,x"0000" -- 68A6
           ,x"0000" -- 68A8
           ,x"0000" -- 68AA
           ,x"0000" -- 68AC
           ,x"0000" -- 68AE
           ,x"0000" -- 68B0
           ,x"0000" -- 68B2
           ,x"0000" -- 68B4
           ,x"0000" -- 68B6
           ,x"0000" -- 68B8
           ,x"0000" -- 68BA
           ,x"0000" -- 68BC
           ,x"0000" -- 68BE
           ,x"0000" -- 68C0
           ,x"0000" -- 68C2
           ,x"0000" -- 68C4
           ,x"0000" -- 68C6
           ,x"0000" -- 68C8
           ,x"0000" -- 68CA
           ,x"0000" -- 68CC
           ,x"0000" -- 68CE
           ,x"0000" -- 68D0
           ,x"0000" -- 68D2
           ,x"0000" -- 68D4
           ,x"0000" -- 68D6
           ,x"0000" -- 68D8
           ,x"0000" -- 68DA
           ,x"0000" -- 68DC
           ,x"0000" -- 68DE
           ,x"0000" -- 68E0
           ,x"0000" -- 68E2
           ,x"0000" -- 68E4
           ,x"0000" -- 68E6
           ,x"0000" -- 68E8
           ,x"0000" -- 68EA
           ,x"0000" -- 68EC
           ,x"0000" -- 68EE
           ,x"0000" -- 68F0
           ,x"0000" -- 68F2
           ,x"0000" -- 68F4
           ,x"0000" -- 68F6
           ,x"0000" -- 68F8
           ,x"0000" -- 68FA
           ,x"0000" -- 68FC
           ,x"0000" -- 68FE
           ,x"0000" -- 6900
           ,x"0000" -- 6902
           ,x"0000" -- 6904
           ,x"0000" -- 6906
           ,x"0000" -- 6908
           ,x"0000" -- 690A
           ,x"0000" -- 690C
           ,x"0000" -- 690E
           ,x"0000" -- 6910
           ,x"0000" -- 6912
           ,x"0000" -- 6914
           ,x"0000" -- 6916
           ,x"0000" -- 6918
           ,x"0000" -- 691A
           ,x"0000" -- 691C
           ,x"0000" -- 691E
           ,x"0000" -- 6920
           ,x"0000" -- 6922
           ,x"0000" -- 6924
           ,x"0000" -- 6926
           ,x"0000" -- 6928
           ,x"0000" -- 692A
           ,x"0000" -- 692C
           ,x"0000" -- 692E
           ,x"0000" -- 6930
           ,x"0000" -- 6932
           ,x"0000" -- 6934
           ,x"0000" -- 6936
           ,x"0000" -- 6938
           ,x"0000" -- 693A
           ,x"0000" -- 693C
           ,x"0000" -- 693E
           ,x"0000" -- 6940
           ,x"0000" -- 6942
           ,x"0000" -- 6944
           ,x"0000" -- 6946
           ,x"0000" -- 6948
           ,x"0000" -- 694A
           ,x"0000" -- 694C
           ,x"0000" -- 694E
           ,x"0000" -- 6950
           ,x"0000" -- 6952
           ,x"0000" -- 6954
           ,x"0000" -- 6956
           ,x"0000" -- 6958
           ,x"0000" -- 695A
           ,x"0000" -- 695C
           ,x"0000" -- 695E
           ,x"0000" -- 6960
           ,x"0000" -- 6962
           ,x"0000" -- 6964
           ,x"0000" -- 6966
           ,x"0000" -- 6968
           ,x"0000" -- 696A
           ,x"0000" -- 696C
           ,x"0000" -- 696E
           ,x"0000" -- 6970
           ,x"0000" -- 6972
           ,x"0000" -- 6974
           ,x"0000" -- 6976
           ,x"0000" -- 6978
           ,x"0000" -- 697A
           ,x"0000" -- 697C
           ,x"0000" -- 697E
           ,x"0000" -- 6980
           ,x"0000" -- 6982
           ,x"0000" -- 6984
           ,x"0000" -- 6986
           ,x"0000" -- 6988
           ,x"0000" -- 698A
           ,x"0000" -- 698C
           ,x"0000" -- 698E
           ,x"0000" -- 6990
           ,x"0000" -- 6992
           ,x"0000" -- 6994
           ,x"0000" -- 6996
           ,x"0000" -- 6998
           ,x"0000" -- 699A
           ,x"0000" -- 699C
           ,x"0000" -- 699E
           ,x"0000" -- 69A0
           ,x"0000" -- 69A2
           ,x"0000" -- 69A4
           ,x"0000" -- 69A6
           ,x"0000" -- 69A8
           ,x"0000" -- 69AA
           ,x"0000" -- 69AC
           ,x"0000" -- 69AE
           ,x"0000" -- 69B0
           ,x"0000" -- 69B2
           ,x"0000" -- 69B4
           ,x"0000" -- 69B6
           ,x"0000" -- 69B8
           ,x"0000" -- 69BA
           ,x"0000" -- 69BC
           ,x"0000" -- 69BE
           ,x"0000" -- 69C0
           ,x"0000" -- 69C2
           ,x"0000" -- 69C4
           ,x"0000" -- 69C6
           ,x"0000" -- 69C8
           ,x"0000" -- 69CA
           ,x"0000" -- 69CC
           ,x"0000" -- 69CE
           ,x"0000" -- 69D0
           ,x"0000" -- 69D2
           ,x"0000" -- 69D4
           ,x"0000" -- 69D6
           ,x"0000" -- 69D8
           ,x"0000" -- 69DA
           ,x"0000" -- 69DC
           ,x"0000" -- 69DE
           ,x"0000" -- 69E0
           ,x"0000" -- 69E2
           ,x"0000" -- 69E4
           ,x"0000" -- 69E6
           ,x"0000" -- 69E8
           ,x"0000" -- 69EA
           ,x"0000" -- 69EC
           ,x"0000" -- 69EE
           ,x"0000" -- 69F0
           ,x"0000" -- 69F2
           ,x"0000" -- 69F4
           ,x"0000" -- 69F6
           ,x"0000" -- 69F8
           ,x"0000" -- 69FA
           ,x"0000" -- 69FC
           ,x"0000" -- 69FE
           ,x"0000" -- 6A00
           ,x"0000" -- 6A02
           ,x"0000" -- 6A04
           ,x"0000" -- 6A06
           ,x"0000" -- 6A08
           ,x"0000" -- 6A0A
           ,x"0000" -- 6A0C
           ,x"0000" -- 6A0E
           ,x"0000" -- 6A10
           ,x"0000" -- 6A12
           ,x"0000" -- 6A14
           ,x"0000" -- 6A16
           ,x"0000" -- 6A18
           ,x"0000" -- 6A1A
           ,x"0000" -- 6A1C
           ,x"0000" -- 6A1E
           ,x"0000" -- 6A20
           ,x"0000" -- 6A22
           ,x"0000" -- 6A24
           ,x"0000" -- 6A26
           ,x"0000" -- 6A28
           ,x"0000" -- 6A2A
           ,x"0000" -- 6A2C
           ,x"0000" -- 6A2E
           ,x"0000" -- 6A30
           ,x"0000" -- 6A32
           ,x"0000" -- 6A34
           ,x"0000" -- 6A36
           ,x"0000" -- 6A38
           ,x"0000" -- 6A3A
           ,x"0000" -- 6A3C
           ,x"0000" -- 6A3E
           ,x"0000" -- 6A40
           ,x"0000" -- 6A42
           ,x"0000" -- 6A44
           ,x"0000" -- 6A46
           ,x"0000" -- 6A48
           ,x"0000" -- 6A4A
           ,x"0000" -- 6A4C
           ,x"0000" -- 6A4E
           ,x"0000" -- 6A50
           ,x"0000" -- 6A52
           ,x"0000" -- 6A54
           ,x"0000" -- 6A56
           ,x"0000" -- 6A58
           ,x"0000" -- 6A5A
           ,x"0000" -- 6A5C
           ,x"0000" -- 6A5E
           ,x"0000" -- 6A60
           ,x"0000" -- 6A62
           ,x"0000" -- 6A64
           ,x"0000" -- 6A66
           ,x"0000" -- 6A68
           ,x"0000" -- 6A6A
           ,x"0000" -- 6A6C
           ,x"0000" -- 6A6E
           ,x"0000" -- 6A70
           ,x"0000" -- 6A72
           ,x"0000" -- 6A74
           ,x"0000" -- 6A76
           ,x"0000" -- 6A78
           ,x"0000" -- 6A7A
           ,x"0000" -- 6A7C
           ,x"0000" -- 6A7E
           ,x"0000" -- 6A80
           ,x"0000" -- 6A82
           ,x"0000" -- 6A84
           ,x"0000" -- 6A86
           ,x"0000" -- 6A88
           ,x"0000" -- 6A8A
           ,x"0000" -- 6A8C
           ,x"0000" -- 6A8E
           ,x"0000" -- 6A90
           ,x"0000" -- 6A92
           ,x"0000" -- 6A94
           ,x"0000" -- 6A96
           ,x"0000" -- 6A98
           ,x"0000" -- 6A9A
           ,x"0000" -- 6A9C
           ,x"0000" -- 6A9E
           ,x"0000" -- 6AA0
           ,x"0000" -- 6AA2
           ,x"0000" -- 6AA4
           ,x"0000" -- 6AA6
           ,x"0000" -- 6AA8
           ,x"0000" -- 6AAA
           ,x"0000" -- 6AAC
           ,x"0000" -- 6AAE
           ,x"0000" -- 6AB0
           ,x"0000" -- 6AB2
           ,x"0000" -- 6AB4
           ,x"0000" -- 6AB6
           ,x"0000" -- 6AB8
           ,x"0000" -- 6ABA
           ,x"0000" -- 6ABC
           ,x"0000" -- 6ABE
           ,x"0000" -- 6AC0
           ,x"0000" -- 6AC2
           ,x"0000" -- 6AC4
           ,x"0000" -- 6AC6
           ,x"0000" -- 6AC8
           ,x"0000" -- 6ACA
           ,x"0000" -- 6ACC
           ,x"0000" -- 6ACE
           ,x"0000" -- 6AD0
           ,x"0000" -- 6AD2
           ,x"0000" -- 6AD4
           ,x"0000" -- 6AD6
           ,x"0000" -- 6AD8
           ,x"0000" -- 6ADA
           ,x"0000" -- 6ADC
           ,x"0000" -- 6ADE
           ,x"0000" -- 6AE0
           ,x"0000" -- 6AE2
           ,x"0000" -- 6AE4
           ,x"0000" -- 6AE6
           ,x"0000" -- 6AE8
           ,x"0000" -- 6AEA
           ,x"0000" -- 6AEC
           ,x"0000" -- 6AEE
           ,x"0000" -- 6AF0
           ,x"0000" -- 6AF2
           ,x"0000" -- 6AF4
           ,x"0000" -- 6AF6
           ,x"0000" -- 6AF8
           ,x"0000" -- 6AFA
           ,x"0000" -- 6AFC
           ,x"0000" -- 6AFE
           ,x"0000" -- 6B00
           ,x"0000" -- 6B02
           ,x"0000" -- 6B04
           ,x"0000" -- 6B06
           ,x"0000" -- 6B08
           ,x"0000" -- 6B0A
           ,x"0000" -- 6B0C
           ,x"0000" -- 6B0E
           ,x"0000" -- 6B10
           ,x"0000" -- 6B12
           ,x"0000" -- 6B14
           ,x"0000" -- 6B16
           ,x"0000" -- 6B18
           ,x"0000" -- 6B1A
           ,x"0000" -- 6B1C
           ,x"0000" -- 6B1E
           ,x"0000" -- 6B20
           ,x"0000" -- 6B22
           ,x"0000" -- 6B24
           ,x"0000" -- 6B26
           ,x"0000" -- 6B28
           ,x"0000" -- 6B2A
           ,x"0000" -- 6B2C
           ,x"0000" -- 6B2E
           ,x"0000" -- 6B30
           ,x"0000" -- 6B32
           ,x"0000" -- 6B34
           ,x"0000" -- 6B36
           ,x"0000" -- 6B38
           ,x"0000" -- 6B3A
           ,x"0000" -- 6B3C
           ,x"0000" -- 6B3E
           ,x"0000" -- 6B40
           ,x"0000" -- 6B42
           ,x"0000" -- 6B44
           ,x"0000" -- 6B46
           ,x"0000" -- 6B48
           ,x"0000" -- 6B4A
           ,x"0000" -- 6B4C
           ,x"0000" -- 6B4E
           ,x"0000" -- 6B50
           ,x"0000" -- 6B52
           ,x"0000" -- 6B54
           ,x"0000" -- 6B56
           ,x"0000" -- 6B58
           ,x"0000" -- 6B5A
           ,x"0000" -- 6B5C
           ,x"0000" -- 6B5E
           ,x"0000" -- 6B60
           ,x"0000" -- 6B62
           ,x"0000" -- 6B64
           ,x"0000" -- 6B66
           ,x"0000" -- 6B68
           ,x"0000" -- 6B6A
           ,x"0000" -- 6B6C
           ,x"0000" -- 6B6E
           ,x"0000" -- 6B70
           ,x"0000" -- 6B72
           ,x"0000" -- 6B74
           ,x"0000" -- 6B76
           ,x"0000" -- 6B78
           ,x"0000" -- 6B7A
           ,x"0000" -- 6B7C
           ,x"0000" -- 6B7E
           ,x"0000" -- 6B80
           ,x"0000" -- 6B82
           ,x"0000" -- 6B84
           ,x"0000" -- 6B86
           ,x"0000" -- 6B88
           ,x"0000" -- 6B8A
           ,x"0000" -- 6B8C
           ,x"0000" -- 6B8E
           ,x"0000" -- 6B90
           ,x"0000" -- 6B92
           ,x"0000" -- 6B94
           ,x"0000" -- 6B96
           ,x"0000" -- 6B98
           ,x"0000" -- 6B9A
           ,x"0000" -- 6B9C
           ,x"0000" -- 6B9E
           ,x"0000" -- 6BA0
           ,x"0000" -- 6BA2
           ,x"0000" -- 6BA4
           ,x"0000" -- 6BA6
           ,x"0000" -- 6BA8
           ,x"0000" -- 6BAA
           ,x"0000" -- 6BAC
           ,x"0000" -- 6BAE
           ,x"0000" -- 6BB0
           ,x"0000" -- 6BB2
           ,x"0000" -- 6BB4
           ,x"0000" -- 6BB6
           ,x"0000" -- 6BB8
           ,x"0000" -- 6BBA
           ,x"0000" -- 6BBC
           ,x"0000" -- 6BBE
           ,x"0000" -- 6BC0
           ,x"0000" -- 6BC2
           ,x"0000" -- 6BC4
           ,x"0000" -- 6BC6
           ,x"0000" -- 6BC8
           ,x"0000" -- 6BCA
           ,x"0000" -- 6BCC
           ,x"0000" -- 6BCE
           ,x"0000" -- 6BD0
           ,x"0000" -- 6BD2
           ,x"0000" -- 6BD4
           ,x"0000" -- 6BD6
           ,x"0000" -- 6BD8
           ,x"0000" -- 6BDA
           ,x"0000" -- 6BDC
           ,x"0000" -- 6BDE
           ,x"0000" -- 6BE0
           ,x"0000" -- 6BE2
           ,x"0000" -- 6BE4
           ,x"0000" -- 6BE6
           ,x"0000" -- 6BE8
           ,x"0000" -- 6BEA
           ,x"0000" -- 6BEC
           ,x"0000" -- 6BEE
           ,x"0000" -- 6BF0
           ,x"0000" -- 6BF2
           ,x"0000" -- 6BF4
           ,x"0000" -- 6BF6
           ,x"0000" -- 6BF8
           ,x"0000" -- 6BFA
           ,x"0000" -- 6BFC
           ,x"0000" -- 6BFE
           ,x"0000" -- 6C00
           ,x"0000" -- 6C02
           ,x"0000" -- 6C04
           ,x"0000" -- 6C06
           ,x"0000" -- 6C08
           ,x"0000" -- 6C0A
           ,x"0000" -- 6C0C
           ,x"0000" -- 6C0E
           ,x"0000" -- 6C10
           ,x"0000" -- 6C12
           ,x"0000" -- 6C14
           ,x"0000" -- 6C16
           ,x"0000" -- 6C18
           ,x"0000" -- 6C1A
           ,x"0000" -- 6C1C
           ,x"0000" -- 6C1E
           ,x"0000" -- 6C20
           ,x"0000" -- 6C22
           ,x"0000" -- 6C24
           ,x"0000" -- 6C26
           ,x"0000" -- 6C28
           ,x"0000" -- 6C2A
           ,x"0000" -- 6C2C
           ,x"0000" -- 6C2E
           ,x"0000" -- 6C30
           ,x"0000" -- 6C32
           ,x"0000" -- 6C34
           ,x"0000" -- 6C36
           ,x"0000" -- 6C38
           ,x"0000" -- 6C3A
           ,x"0000" -- 6C3C
           ,x"0000" -- 6C3E
           ,x"0000" -- 6C40
           ,x"0000" -- 6C42
           ,x"0000" -- 6C44
           ,x"0000" -- 6C46
           ,x"0000" -- 6C48
           ,x"0000" -- 6C4A
           ,x"0000" -- 6C4C
           ,x"0000" -- 6C4E
           ,x"0000" -- 6C50
           ,x"0000" -- 6C52
           ,x"0000" -- 6C54
           ,x"0000" -- 6C56
           ,x"0000" -- 6C58
           ,x"0000" -- 6C5A
           ,x"0000" -- 6C5C
           ,x"0000" -- 6C5E
           ,x"0000" -- 6C60
           ,x"0000" -- 6C62
           ,x"0000" -- 6C64
           ,x"0000" -- 6C66
           ,x"0000" -- 6C68
           ,x"0000" -- 6C6A
           ,x"0000" -- 6C6C
           ,x"0000" -- 6C6E
           ,x"0000" -- 6C70
           ,x"0000" -- 6C72
           ,x"0000" -- 6C74
           ,x"0000" -- 6C76
           ,x"0000" -- 6C78
           ,x"0000" -- 6C7A
           ,x"0000" -- 6C7C
           ,x"0000" -- 6C7E
           ,x"0000" -- 6C80
           ,x"0000" -- 6C82
           ,x"0000" -- 6C84
           ,x"0000" -- 6C86
           ,x"0000" -- 6C88
           ,x"0000" -- 6C8A
           ,x"0000" -- 6C8C
           ,x"0000" -- 6C8E
           ,x"0000" -- 6C90
           ,x"0000" -- 6C92
           ,x"0000" -- 6C94
           ,x"0000" -- 6C96
           ,x"0000" -- 6C98
           ,x"0000" -- 6C9A
           ,x"0000" -- 6C9C
           ,x"0000" -- 6C9E
           ,x"0000" -- 6CA0
           ,x"0000" -- 6CA2
           ,x"0000" -- 6CA4
           ,x"0000" -- 6CA6
           ,x"0000" -- 6CA8
           ,x"0000" -- 6CAA
           ,x"0000" -- 6CAC
           ,x"0000" -- 6CAE
           ,x"0000" -- 6CB0
           ,x"0000" -- 6CB2
           ,x"0000" -- 6CB4
           ,x"0000" -- 6CB6
           ,x"0000" -- 6CB8
           ,x"934b" -- 6CBA
           ,x"2449" -- 6CBC
           ,x"2300" -- 6CBE
           ,x"6204" -- 6CC0
           ,x"08e8" -- 6CC2
           ,x"e280" -- 6CC4
           ,x"6204" -- 6CC6
           ,x"08e8" -- 6CC8
           ,x"4280" -- 6CCA
           ,x"e20e" -- 6CCC
           ,x"20e8" -- 6CCE
           ,x"e280" -- 6CD0
           ,x"e20e" -- 6CD2
           ,x"20e8" -- 6CD4
           ,x"4100" -- 6CD6
           ,x"e20d" -- 6CD8
           ,x"2ae8" -- 6CDA
           ,x"a180" -- 6CDC
           ,x"624f" -- 6CDE
           ,x"2428" -- 6CE0
           ,x"c280" -- 6CE2
           ,x"628c" -- 6CE4
           ,x"28d0" -- 6CE6
           ,x"4180" -- 6CE8
           ,x"628d" -- 6CEA
           ,x"a8d0" -- 6CEC
           ,x"2300" -- 6CEE
           ,x"a38a" -- 6CF0
           ,x"0038" -- 6CF2
           ,x"4100" -- 6CF4
           ,x"820b" -- 6CF6
           ,x"a8f0" -- 6CF8
           ,x"8200" -- 6CFA
           ,x"8942" -- 6CFC
           ,x"0038" -- 6CFE
           ,x"4100" -- 6D00
           ,x"e20f" -- 6D02
           ,x"a8b0" -- 6D04
           ,x"8200" -- 6D06
           ,x"6208" -- 6D08
           ,x"1c49" -- 6D0A
           ,x"c480" -- 6D0C
           ,x"6205" -- 6D0E
           ,x"0ae8" -- 6D10
           ,x"a100" -- 6D12
           ,x"6204" -- 6D14
           ,x"0ed0" -- 6D16
           ,x"4380" -- 6D18
           ,x"c28a" -- 6D1A
           ,x"3020" -- 6D1C
           ,x"8380" -- 6D1E
           ,x"c28a" -- 6D20
           ,x"3010" -- 6D22
           ,x"4100" -- 6D24
           ,x"c28b" -- 6D26
           ,x"3210" -- 6D28
           ,x"8380" -- 6D2A
           ,x"c28b" -- 6D2C
           ,x"3210" -- 6D2E
           ,x"2300" -- 6D30
           ,x"c28a" -- 6D32
           ,x"3218" -- 6D34
           ,x"e080" -- 6D36
           ,x"d2c9" -- 6D38
           ,x"0828" -- 6D3A
           ,x"c280" -- 6D3C
           ,x"6204" -- 6D3E
           ,x"0ad0" -- 6D40
           ,x"4100" -- 6D42
           ,x"e20f" -- 6D44
           ,x"2af0" -- 6D46
           ,x"a300" -- 6D48
           ,x"6206" -- 6D4A
           ,x"1269" -- 6D4C
           ,x"6480" -- 6D4E
           ,x"e20e" -- 6D50
           ,x"20eb" -- 6D52
           ,x"6a80" -- 6D54
           ,x"6207" -- 6D56
           ,x"0af0" -- 6D58
           ,x"a300" -- 6D5A
           ,x"e20e" -- 6D5C
           ,x"26e0" -- 6D5E
           ,x"8180" -- 6D60
           ,x"e20d" -- 6D62
           ,x"a890" -- 6D64
           ,x"2300" -- 6D66
           ,x"6209" -- 6D68
           ,x"ac91" -- 6D6A
           ,x"a300" -- 6D6C
           ,x"e28d" -- 6D6E
           ,x"a810" -- 6D70
           ,x"2300" -- 6D72
           ,x"a28b" -- 6D74
           ,x"9810" -- 6D76
           ,x"2300" -- 6D78
           ,x"0000" -- 6D7A
           ,x"0000" -- 6D7C
           ,x"0000" -- 6D7E
           ,x"2082" -- 6D80
           ,x"0820" -- 6D82
           ,x"0200" -- 6D84
           ,x"5145" -- 6D86
           ,x"0000" -- 6D88
           ,x"0000" -- 6D8A
           ,x"514f" -- 6D8C
           ,x"94f9" -- 6D8E
           ,x"4500" -- 6D90
           ,x"21ea" -- 6D92
           ,x"1c2b" -- 6D94
           ,x"c200" -- 6D96
           ,x"c321" -- 6D98
           ,x"0842" -- 6D9A
           ,x"6180" -- 6D9C
           ,x"428a" -- 6D9E
           ,x"10aa" -- 6DA0
           ,x"4680" -- 6DA2
           ,x"1084" -- 6DA4
           ,x"0000" -- 6DA6
           ,x"0000" -- 6DA8
           ,x"2108" -- 6DAA
           ,x"2081" -- 6DAC
           ,x"0200" -- 6DAE
           ,x"2040" -- 6DB0
           ,x"8208" -- 6DB2
           ,x"4200" -- 6DB4
           ,x"22a7" -- 6DB6
           ,x"3e72" -- 6DB8
           ,x"a200" -- 6DBA
           ,x"0082" -- 6DBC
           ,x"3e20" -- 6DBE
           ,x"8000" -- 6DC0
           ,x"0000" -- 6DC2
           ,x"0020" -- 6DC4
           ,x"8400" -- 6DC6
           ,x"0000" -- 6DC8
           ,x"3e00" -- 6DCA
           ,x"0000" -- 6DCC
           ,x"0000" -- 6DCE
           ,x"0000" -- 6DD0
           ,x"0200" -- 6DD2
           ,x"0021" -- 6DD4
           ,x"0842" -- 6DD6
           ,x"0000" -- 6DD8
           ,x"7229" -- 6DDA
           ,x"aaca" -- 6DDC
           ,x"2700" -- 6DDE
           ,x"2182" -- 6DE0
           ,x"0820" -- 6DE2
           ,x"8700" -- 6DE4
           ,x"7220" -- 6DE6
           ,x"8c42" -- 6DE8
           ,x"0f80" -- 6DEA
           ,x"7220" -- 6DEC
           ,x"8c0a" -- 6DEE
           ,x"2700" -- 6DF0
           ,x"10c5" -- 6DF2
           ,x"24f8" -- 6DF4
           ,x"4100" -- 6DF6
           ,x"fa0f" -- 6DF8
           ,x"020a" -- 6DFA
           ,x"2700" -- 6DFC
           ,x"3908" -- 6DFE
           ,x"3c8a" -- 6E00
           ,x"2700" -- 6E02
           ,x"f821" -- 6E04
           ,x"0841" -- 6E06
           ,x"0400" -- 6E08
           ,x"7228" -- 6E0A
           ,x"9c8a" -- 6E0C
           ,x"2700" -- 6E0E
           ,x"7228" -- 6E10
           ,x"9e08" -- 6E12
           ,x"4e00" -- 6E14
           ,x"0002" -- 6E16
           ,x"0020" -- 6E18
           ,x"0000" -- 6E1A
           ,x"0002" -- 6E1C
           ,x"0020" -- 6E1E
           ,x"8400" -- 6E20
           ,x"1084" -- 6E22
           ,x"2040" -- 6E24
           ,x"8100" -- 6E26
           ,x"000f" -- 6E28
           ,x"80f8" -- 6E2A
           ,x"0000" -- 6E2C
           ,x"4081" -- 6E2E
           ,x"0210" -- 6E30
           ,x"8400" -- 6E32
           ,x"7221" -- 6E34
           ,x"0820" -- 6E36
           ,x"0200" -- 6E38
           ,x"722b" -- 6E3A
           ,x"aaba" -- 6E3C
           ,x"0780" -- 6E3E
           ,x"7228" -- 6E40
           ,x"be8a" -- 6E42
           ,x"2880" -- 6E44
           ,x"f124" -- 6E46
           ,x"9c49" -- 6E48
           ,x"2f00" -- 6E4A
           ,x"7228" -- 6E4C
           ,x"2082" -- 6E4E
           ,x"2700" -- 6E50
           ,x"f124" -- 6E52
           ,x"9249" -- 6E54
           ,x"2f00" -- 6E56
           ,x"fa08" -- 6E58
           ,x"3c82" -- 6E5A
           ,x"0f80" -- 6E5C
           ,x"fa08" -- 6E5E
           ,x"3c82" -- 6E60
           ,x"0800" -- 6E62
           ,x"7a08" -- 6E64
           ,x"209a" -- 6E66
           ,x"2780" -- 6E68
           ,x"8a28" -- 6E6A
           ,x"be8a" -- 6E6C
           ,x"2880" -- 6E6E
           ,x"7082" -- 6E70
           ,x"0820" -- 6E72
           ,x"8700" -- 6E74
           ,x"0820" -- 6E76
           ,x"820a" -- 6E78
           ,x"2700" -- 6E7A
           ,x"8a4a" -- 6E7C
           ,x"30a2" -- 6E7E
           ,x"4880" -- 6E80
           ,x"8208" -- 6E82
           ,x"2082" -- 6E84
           ,x"0f80" -- 6E86
           ,x"8b6a" -- 6E88
           ,x"aa8a" -- 6E8A
           ,x"2880" -- 6E8C
           ,x"8a2c" -- 6E8E
           ,x"aa9a" -- 6E90
           ,x"2880" -- 6E92
           ,x"fa28" -- 6E94
           ,x"a28a" -- 6E96
           ,x"2f80" -- 6E98
           ,x"f228" -- 6E9A
           ,x"bc82" -- 6E9C
           ,x"0800" -- 6E9E
           ,x"7228" -- 6EA0
           ,x"a2aa" -- 6EA2
           ,x"4680" -- 6EA4
           ,x"f228" -- 6EA6
           ,x"bca2" -- 6EA8
           ,x"4880" -- 6EAA
           ,x"7228" -- 6EAC
           ,x"1c0a" -- 6EAE
           ,x"2700" -- 6EB0
           ,x"f882" -- 6EB2
           ,x"0820" -- 6EB4
           ,x"8200" -- 6EB6
           ,x"8a28" -- 6EB8
           ,x"a28a" -- 6EBA
           ,x"2700" -- 6EBC
           ,x"8a28" -- 6EBE
           ,x"9450" -- 6EC0
           ,x"8200" -- 6EC2
           ,x"8a28" -- 6EC4
           ,x"aaaa" -- 6EC6
           ,x"a500" -- 6EC8
           ,x"8a25" -- 6ECA
           ,x"0852" -- 6ECC
           ,x"2880" -- 6ECE
           ,x"8a25" -- 6ED0
           ,x"0820" -- 6ED2
           ,x"8200" -- 6ED4
           ,x"f821" -- 6ED6
           ,x"0842" -- 6ED8
           ,x"0f80" -- 6EDA
           ,x"3882" -- 6EDC
           ,x"0820" -- 6EDE
           ,x"8380" -- 6EE0
           ,x"0204" -- 6EE2
           ,x"0810" -- 6EE4
           ,x"2000" -- 6EE6
           ,x"7041" -- 6EE8
           ,x"0410" -- 6EEA
           ,x"4700" -- 6EEC
           ,x"2148" -- 6EEE
           ,x"8000" -- 6EF0
           ,x"0000" -- 6EF2
           ,x"0000" -- 6EF4
           ,x"0000" -- 6EF6
           ,x"0f80" -- 6EF8
           ,x"4081" -- 6EFA
           ,x"0000" -- 6EFC
           ,x"0000" -- 6EFE
           ,x"0007" -- 6F00
           ,x"22fa" -- 6F02
           ,x"2880" -- 6F04
           ,x"000f" -- 6F06
           ,x"1271" -- 6F08
           ,x"2f00" -- 6F0A
           ,x"0007" -- 6F0C
           ,x"a082" -- 6F0E
           ,x"0780" -- 6F10
           ,x"000f" -- 6F12
           ,x"1249" -- 6F14
           ,x"2f00" -- 6F16
           ,x"000f" -- 6F18
           ,x"20e2" -- 6F1A
           ,x"0f00" -- 6F1C
           ,x"000f" -- 6F1E
           ,x"20e2" -- 6F20
           ,x"0800" -- 6F22
           ,x"0007" -- 6F24
           ,x"a0ba" -- 6F26
           ,x"2700" -- 6F28
           ,x"0008" -- 6F2A
           ,x"a2fa" -- 6F2C
           ,x"2880" -- 6F2E
           ,x"0007" -- 6F30
           ,x"0820" -- 6F32
           ,x"8700" -- 6F34
           ,x"0007" -- 6F36
           ,x"0822" -- 6F38
           ,x"8e00" -- 6F3A
           ,x"0009" -- 6F3C
           ,x"28c2" -- 6F3E
           ,x"8900" -- 6F40
           ,x"0008" -- 6F42
           ,x"2082" -- 6F44
           ,x"0f80" -- 6F46
           ,x"0008" -- 6F48
           ,x"b6aa" -- 6F4A
           ,x"2880" -- 6F4C
           ,x"0008" -- 6F4E
           ,x"b2aa" -- 6F50
           ,x"6880" -- 6F52
           ,x"000f" -- 6F54
           ,x"a28a" -- 6F56
           ,x"2f80" -- 6F58
           ,x"000f" -- 6F5A
           ,x"22f2" -- 6F5C
           ,x"0800" -- 6F5E
           ,x"000f" -- 6F60
           ,x"a2aa" -- 6F62
           ,x"4e80" -- 6F64
           ,x"000f" -- 6F66
           ,x"22f2" -- 6F68
           ,x"8900" -- 6F6A
           ,x"0007" -- 6F6C
           ,x"a070" -- 6F6E
           ,x"2f00" -- 6F70
           ,x"000f" -- 6F72
           ,x"8820" -- 6F74
           ,x"8200" -- 6F76
           ,x"0004" -- 6F78
           ,x"9249" -- 6F7A
           ,x"2300" -- 6F7C
           ,x"0008" -- 6F7E
           ,x"a292" -- 6F80
           ,x"8400" -- 6F82
           ,x"0008" -- 6F84
           ,x"a2ab" -- 6F86
           ,x"6880" -- 6F88
           ,x"0008" -- 6F8A
           ,x"9421" -- 6F8C
           ,x"4880" -- 6F8E
           ,x"0008" -- 6F90
           ,x"9420" -- 6F92
           ,x"8200" -- 6F94
           ,x"000f" -- 6F96
           ,x"8421" -- 6F98
           ,x"0f80" -- 6F9A
           ,x"3104" -- 6F9C
           ,x"2041" -- 6F9E
           ,x"0300" -- 6FA0
           ,x"2082" -- 6FA2
           ,x"0020" -- 6FA4
           ,x"8200" -- 6FA6
           ,x"6041" -- 6FA8
           ,x"0210" -- 6FAA
           ,x"4600" -- 6FAC
           ,x"42a1" -- 6FAE
           ,x"0000" -- 6FB0
           ,x"0000" -- 6FB2
           ,x"8ddb" -- 6FB4
           ,x"f7df" -- 6FB6
           ,x"fdff" -- 6FB8
           ,x"0000" -- 6FBA
           ,x"0000" -- 6FBC
           ,x"001c" -- 6FBE
           ,x"0000" -- 6FC0
           ,x"0000" -- 6FC2
           ,x"071c" -- 6FC4
           ,x"0000" -- 6FC6
           ,x"0001" -- 6FC8
           ,x"c71c" -- 6FCA
           ,x"0000" -- 6FCC
           ,x"0071" -- 6FCE
           ,x"c71c" -- 6FD0
           ,x"0000" -- 6FD2
           ,x"1c71" -- 6FD4
           ,x"c71c" -- 6FD6
           ,x"0007" -- 6FD8
           ,x"1c71" -- 6FDA
           ,x"c71c" -- 6FDC
           ,x"01c7" -- 6FDE
           ,x"1c71" -- 6FE0
           ,x"c71c" -- 6FE2
           ,x"71c7" -- 6FE4
           ,x"1c71" -- 6FE6
           ,x"c71c" -- 6FE8
           ,x"7a1b" -- 6FEA
           ,x"69b6" -- 6FEC
           ,x"1780" -- 6FEE
           ,x"a95a" -- 6FF0
           ,x"95a9" -- 6FF2
           ,x"5a95" -- 6FF4
           ,x"0007" -- 6FF6
           ,x"df7d" -- 6FF8
           ,x"c71c" -- 6FFA
           ,x"71cf" -- 6FFC
           ,x"3cf1" -- 6FFE
           ,x"c71c" -- 7000
           ,x"000f" -- 7002
           ,x"fffd" -- 7004
           ,x"c71c" -- 7006
           ,x"71c7" -- 7008
           ,x"df7c" -- 700A
           ,x"0000" -- 700C
           ,x"0c61" -- 700E
           ,x"0821" -- 7010
           ,x"0c20" -- 7012
           ,x"03f0" -- 7014
           ,x"0003" -- 7016
           ,x"f000" -- 7018
           ,x"0008" -- 701A
           ,x"2080" -- 701C
           ,x"0000" -- 701E
           ,x"000c" -- 7020
           ,x"30c0" -- 7022
           ,x"0000" -- 7024
           ,x"000e" -- 7026
           ,x"38e0" -- 7028
           ,x"0000" -- 702A
           ,x"000f" -- 702C
           ,x"3cf0" -- 702E
           ,x"0000" -- 7030
           ,x"000f" -- 7032
           ,x"bef8" -- 7034
           ,x"0000" -- 7036
           ,x"000f" -- 7038
           ,x"fffc" -- 703A
           ,x"0000" -- 703C
           ,x"3124" -- 703E
           ,x"1c41" -- 7040
           ,x"0b80" -- 7042
           ,x"0007" -- 7044
           ,x"1c70" -- 7046
           ,x"0000" -- 7048
           ,x"71cf" -- 704A
           ,x"fffd" -- 704C
           ,x"c71c" -- 704E
           ,x"ffff" -- 7050
           ,x"ffff" -- 7052
           ,x"ffff" -- 7054
           ,x"000f" -- 7056
           ,x"3cf1" -- 7058
           ,x"c71c" -- 705A
           ,x"71c7" -- 705C
           ,x"df7d" -- 705E
           ,x"c71c" -- 7060
           ,x"71cf" -- 7062
           ,x"fffc" -- 7064
           ,x"0000" -- 7066
           ,x"71cf" -- 7068
           ,x"3cf0" -- 706A
           ,x"0000" -- 706C
           ,x"8304" -- 706E
           ,x"0820" -- 7070
           ,x"4183" -- 7072
           ,x"8a28" -- 7074
           ,x"a28a" -- 7076
           ,x"28a2" -- 7078
           ,x"21ca" -- 707A
           ,x"8820" -- 707C
           ,x"8200" -- 707E
           ,x"2082" -- 7080
           ,x"08a9" -- 7082
           ,x"c200" -- 7084
           ,x"0081" -- 7086
           ,x"3e10" -- 7088
           ,x"8000" -- 708A
           ,x"0084" -- 708C
           ,x"3e40" -- 708E
           ,x"8000" -- 7090
           ,x"00e1" -- 7092
           ,x"8a42" -- 7094
           ,x"0000" -- 7096
           ,x"0021" -- 7098
           ,x"28c3" -- 709A
           ,x"8000" -- 709C
           ,x"0204" -- 709E
           ,x"0a18" -- 70A0
           ,x"e000" -- 70A2
           ,x"038c" -- 70A4
           ,x"2810" -- 70A6
           ,x"2000" -- 70A8
           ,x"21c2" -- 70AA
           ,x"2aa9" -- 70AC
           ,x"c000" -- 70AE
           ,x"ffff" -- 70B0
           ,x"ffff" -- 70B2
           ,x"ffff" -- 70B4
           ,x"ffff" -- 70B6
           ,x"ffff" -- 70B8
           ,x"ffff" -- 70BA
           ,x"ffff" -- 70BC
           ,x"ffff" -- 70BE
           ,x"ffff" -- 70C0
           ,x"ffff" -- 70C2
           ,x"ffff" -- 70C4
           ,x"ffff" -- 70C6
           ,x"ffff" -- 70C8
           ,x"ffff" -- 70CA
           ,x"ffff" -- 70CC
           ,x"ffff" -- 70CE
           ,x"ffff" -- 70D0
           ,x"ffff" -- 70D2
           ,x"ffff" -- 70D4
           ,x"ffff" -- 70D6
           ,x"ffff" -- 70D8
           ,x"ffff" -- 70DA
           ,x"ffff" -- 70DC
           ,x"ffff" -- 70DE
           ,x"ffff" -- 70E0
           ,x"ffff" -- 70E2
           ,x"ffff" -- 70E4
           ,x"ffff" -- 70E6
           ,x"ffff" -- 70E8
           ,x"ffff" -- 70EA
           ,x"ffff" -- 70EC
           ,x"ffff" -- 70EE
           ,x"ffff" -- 70F0
           ,x"ffff" -- 70F2
           ,x"ffff" -- 70F4
           ,x"ffff" -- 70F6
           ,x"ffff" -- 70F8
           ,x"ffff" -- 70FA
           ,x"ffff" -- 70FC
           ,x"ffff" -- 70FE
           ,x"ffff" -- 7100
           ,x"ffff" -- 7102
           ,x"ffff" -- 7104
           ,x"ffff" -- 7106
           ,x"ffff" -- 7108
           ,x"ffff" -- 710A
           ,x"ffff" -- 710C
           ,x"ffff" -- 710E
           ,x"ffff" -- 7110
           ,x"ffff" -- 7112
           ,x"ffff" -- 7114
           ,x"ffff" -- 7116
           ,x"ffff" -- 7118
           ,x"ffff" -- 711A
           ,x"ffff" -- 711C
           ,x"ffff" -- 711E
           ,x"ffff" -- 7120
           ,x"ffff" -- 7122
           ,x"ffff" -- 7124
           ,x"ffff" -- 7126
           ,x"ffff" -- 7128
           ,x"ffff" -- 712A
           ,x"ffff" -- 712C
           ,x"ffff" -- 712E
           ,x"ffff" -- 7130
           ,x"ffff" -- 7132
           ,x"ffff" -- 7134
           ,x"ffff" -- 7136
           ,x"ffff" -- 7138
           ,x"ffff" -- 713A
           ,x"ffff" -- 713C
           ,x"ffff" -- 713E
           ,x"ffff" -- 7140
           ,x"ffff" -- 7142
           ,x"ffff" -- 7144
           ,x"ffff" -- 7146
           ,x"ffff" -- 7148
           ,x"ffff" -- 714A
           ,x"ffff" -- 714C
           ,x"ffff" -- 714E
           ,x"ffff" -- 7150
           ,x"ffff" -- 7152
           ,x"ffff" -- 7154
           ,x"ffff" -- 7156
           ,x"ffff" -- 7158
           ,x"ffff" -- 715A
           ,x"ffff" -- 715C
           ,x"ffff" -- 715E
           ,x"ffff" -- 7160
           ,x"ffff" -- 7162
           ,x"ffff" -- 7164
           ,x"ffff" -- 7166
           ,x"ffff" -- 7168
           ,x"ffff" -- 716A
           ,x"ffff" -- 716C
           ,x"ffff" -- 716E
           ,x"ffff" -- 7170
           ,x"ffff" -- 7172
           ,x"ffff" -- 7174
           ,x"ffff" -- 7176
           ,x"ffff" -- 7178
           ,x"ffff" -- 717A
           ,x"ffff" -- 717C
           ,x"ffff" -- 717E
           ,x"ffff" -- 7180
           ,x"ffff" -- 7182
           ,x"ffff" -- 7184
           ,x"ffff" -- 7186
           ,x"ffff" -- 7188
           ,x"ffff" -- 718A
           ,x"ffff" -- 718C
           ,x"ffff" -- 718E
           ,x"ffff" -- 7190
           ,x"ffff" -- 7192
           ,x"ffff" -- 7194
           ,x"ffff" -- 7196
           ,x"ffff" -- 7198
           ,x"ffff" -- 719A
           ,x"ffff" -- 719C
           ,x"ffff" -- 719E
           ,x"ffff" -- 71A0
           ,x"ffff" -- 71A2
           ,x"ffff" -- 71A4
           ,x"ffff" -- 71A6
           ,x"ffff" -- 71A8
           ,x"ffff" -- 71AA
           ,x"ffff" -- 71AC
           ,x"ffff" -- 71AE
           ,x"ffff" -- 71B0
           ,x"ffff" -- 71B2
           ,x"ffff" -- 71B4
           ,x"ffff" -- 71B6
           ,x"ffff" -- 71B8
           ,x"ffff" -- 71BA
           ,x"ffff" -- 71BC
           ,x"ffff" -- 71BE
           ,x"ffff" -- 71C0
           ,x"ffff" -- 71C2
           ,x"ffff" -- 71C4
           ,x"ffff" -- 71C6
           ,x"ffff" -- 71C8
           ,x"ffff" -- 71CA
           ,x"ffff" -- 71CC
           ,x"ffff" -- 71CE
           ,x"ffff" -- 71D0
           ,x"ffff" -- 71D2
           ,x"ffff" -- 71D4
           ,x"ffff" -- 71D6
           ,x"ffff" -- 71D8
           ,x"ffff" -- 71DA
           ,x"ffff" -- 71DC
           ,x"ffff" -- 71DE
           ,x"ffff" -- 71E0
           ,x"ffff" -- 71E2
           ,x"ffff" -- 71E4
           ,x"ffff" -- 71E6
           ,x"ffff" -- 71E8
           ,x"ffff" -- 71EA
           ,x"ffff" -- 71EC
           ,x"ffff" -- 71EE
           ,x"ffff" -- 71F0
           ,x"ffff" -- 71F2
           ,x"ffff" -- 71F4
           ,x"ffff" -- 71F6
           ,x"ffff" -- 71F8
           ,x"ffff" -- 71FA
           ,x"ffff" -- 71FC
           ,x"ffff" -- 71FE
           ,x"ffff" -- 7200
           ,x"ffff" -- 7202
           ,x"ffff" -- 7204
           ,x"ffff" -- 7206
           ,x"ffff" -- 7208
           ,x"ffff" -- 720A
           ,x"ffff" -- 720C
           ,x"ffff" -- 720E
           ,x"ffff" -- 7210
           ,x"ffff" -- 7212
           ,x"ffff" -- 7214
           ,x"ffff" -- 7216
           ,x"ffff" -- 7218
           ,x"ffff" -- 721A
           ,x"ffff" -- 721C
           ,x"ffff" -- 721E
           ,x"ffff" -- 7220
           ,x"ffff" -- 7222
           ,x"ffff" -- 7224
           ,x"ffff" -- 7226
           ,x"ffff" -- 7228
           ,x"ffff" -- 722A
           ,x"ffff" -- 722C
           ,x"ffff" -- 722E
           ,x"ffff" -- 7230
           ,x"ffff" -- 7232
           ,x"ffff" -- 7234
           ,x"ffff" -- 7236
           ,x"ffff" -- 7238
           ,x"ffff" -- 723A
           ,x"ffff" -- 723C
           ,x"ffff" -- 723E
           ,x"ffff" -- 7240
           ,x"ffff" -- 7242
           ,x"ffff" -- 7244
           ,x"ffff" -- 7246
           ,x"ffff" -- 7248
           ,x"ffff" -- 724A
           ,x"ffff" -- 724C
           ,x"ffff" -- 724E
           ,x"ffff" -- 7250
           ,x"ffff" -- 7252
           ,x"ffff" -- 7254
           ,x"ffff" -- 7256
           ,x"ffff" -- 7258
           ,x"ffff" -- 725A
           ,x"ffff" -- 725C
           ,x"ffff" -- 725E
           ,x"ffff" -- 7260
           ,x"ffff" -- 7262
           ,x"ffff" -- 7264
           ,x"ffff" -- 7266
           ,x"ffff" -- 7268
           ,x"ffff" -- 726A
           ,x"ffff" -- 726C
           ,x"ffff" -- 726E
           ,x"ffff" -- 7270
           ,x"ffff" -- 7272
           ,x"ffff" -- 7274
           ,x"ffff" -- 7276
           ,x"ffff" -- 7278
           ,x"ffff" -- 727A
           ,x"ffff" -- 727C
           ,x"ffff" -- 727E
           ,x"ffff" -- 7280
           ,x"ffff" -- 7282
           ,x"ffff" -- 7284
           ,x"ffff" -- 7286
           ,x"ffff" -- 7288
           ,x"ffff" -- 728A
           ,x"ffff" -- 728C
           ,x"ffff" -- 728E
           ,x"ffff" -- 7290
           ,x"ffff" -- 7292
           ,x"ffff" -- 7294
           ,x"ffff" -- 7296
           ,x"ffff" -- 7298
           ,x"ffff" -- 729A
           ,x"ffff" -- 729C
           ,x"ffff" -- 729E
           ,x"ffff" -- 72A0
           ,x"ffff" -- 72A2
           ,x"ffff" -- 72A4
           ,x"ffff" -- 72A6
           ,x"ffff" -- 72A8
           ,x"ffff" -- 72AA
           ,x"ffff" -- 72AC
           ,x"ffff" -- 72AE
           ,x"ffff" -- 72B0
           ,x"ffff" -- 72B2
           ,x"ffff" -- 72B4
           ,x"ffff" -- 72B6
           ,x"ffff" -- 72B8
           ,x"ffff" -- 72BA
           ,x"ffff" -- 72BC
           ,x"ffff" -- 72BE
           ,x"ffff" -- 72C0
           ,x"ffff" -- 72C2
           ,x"ffff" -- 72C4
           ,x"ffff" -- 72C6
           ,x"ffff" -- 72C8
           ,x"ffff" -- 72CA
           ,x"ffff" -- 72CC
           ,x"ffff" -- 72CE
           ,x"ffff" -- 72D0
           ,x"ffff" -- 72D2
           ,x"ffff" -- 72D4
           ,x"ffff" -- 72D6
           ,x"ffff" -- 72D8
           ,x"ffff" -- 72DA
           ,x"ffff" -- 72DC
           ,x"ffff" -- 72DE
           ,x"ffff" -- 72E0
           ,x"ffff" -- 72E2
           ,x"ffff" -- 72E4
           ,x"ffff" -- 72E6
           ,x"ffff" -- 72E8
           ,x"ffff" -- 72EA
           ,x"ffff" -- 72EC
           ,x"ffff" -- 72EE
           ,x"ffff" -- 72F0
           ,x"ffff" -- 72F2
           ,x"ffff" -- 72F4
           ,x"ffff" -- 72F6
           ,x"ffff" -- 72F8
           ,x"ffff" -- 72FA
           ,x"ffff" -- 72FC
           ,x"ffff" -- 72FE
           ,x"ffff" -- 7300
           ,x"ffff" -- 7302
           ,x"ffff" -- 7304
           ,x"ffff" -- 7306
           ,x"ffff" -- 7308
           ,x"ffff" -- 730A
           ,x"ffff" -- 730C
           ,x"ffff" -- 730E
           ,x"ffff" -- 7310
           ,x"ffff" -- 7312
           ,x"ffff" -- 7314
           ,x"ffff" -- 7316
           ,x"ffff" -- 7318
           ,x"ffff" -- 731A
           ,x"ffff" -- 731C
           ,x"ffff" -- 731E
           ,x"ffff" -- 7320
           ,x"ffff" -- 7322
           ,x"ffff" -- 7324
           ,x"ffff" -- 7326
           ,x"ffff" -- 7328
           ,x"ffff" -- 732A
           ,x"ffff" -- 732C
           ,x"ffff" -- 732E
           ,x"ffff" -- 7330
           ,x"ffff" -- 7332
           ,x"ffff" -- 7334
           ,x"ffff" -- 7336
           ,x"ffff" -- 7338
           ,x"ffff" -- 733A
           ,x"ffff" -- 733C
           ,x"ffff" -- 733E
           ,x"ffff" -- 7340
           ,x"ffff" -- 7342
           ,x"ffff" -- 7344
           ,x"ffff" -- 7346
           ,x"ffff" -- 7348
           ,x"ffff" -- 734A
           ,x"ffff" -- 734C
           ,x"ffff" -- 734E
           ,x"ffff" -- 7350
           ,x"ffff" -- 7352
           ,x"ffff" -- 7354
           ,x"ffff" -- 7356
           ,x"ffff" -- 7358
           ,x"ffff" -- 735A
           ,x"ffff" -- 735C
           ,x"ffff" -- 735E
           ,x"ffff" -- 7360
           ,x"ffff" -- 7362
           ,x"ffff" -- 7364
           ,x"ffff" -- 7366
           ,x"ffff" -- 7368
           ,x"ffff" -- 736A
           ,x"ffff" -- 736C
           ,x"ffff" -- 736E
           ,x"ffff" -- 7370
           ,x"ffff" -- 7372
           ,x"ffff" -- 7374
           ,x"ffff" -- 7376
           ,x"ffff" -- 7378
           ,x"ffff" -- 737A
           ,x"ffff" -- 737C
           ,x"ffff" -- 737E
           ,x"ffff" -- 7380
           ,x"ffff" -- 7382
           ,x"ffff" -- 7384
           ,x"ffff" -- 7386
           ,x"ffff" -- 7388
           ,x"ffff" -- 738A
           ,x"ffff" -- 738C
           ,x"ffff" -- 738E
           ,x"ffff" -- 7390
           ,x"ffff" -- 7392
           ,x"ffff" -- 7394
           ,x"ffff" -- 7396
           ,x"ffff" -- 7398
           ,x"ffff" -- 739A
           ,x"ffff" -- 739C
           ,x"ffff" -- 739E
           ,x"ffff" -- 73A0
           ,x"ffff" -- 73A2
           ,x"ffff" -- 73A4
           ,x"ffff" -- 73A6
           ,x"ffff" -- 73A8
           ,x"ffff" -- 73AA
           ,x"ffff" -- 73AC
           ,x"ffff" -- 73AE
           ,x"ffff" -- 73B0
           ,x"ffff" -- 73B2
           ,x"ffff" -- 73B4
           ,x"ffff" -- 73B6
           ,x"ffff" -- 73B8
           ,x"ffff" -- 73BA
           ,x"ffff" -- 73BC
           ,x"ffff" -- 73BE
           ,x"ffff" -- 73C0
           ,x"ffff" -- 73C2
           ,x"ffff" -- 73C4
           ,x"ffff" -- 73C6
           ,x"ffff" -- 73C8
           ,x"ffff" -- 73CA
           ,x"ffff" -- 73CC
           ,x"ffff" -- 73CE
           ,x"ffff" -- 73D0
           ,x"ffff" -- 73D2
           ,x"ffff" -- 73D4
           ,x"ffff" -- 73D6
           ,x"ffff" -- 73D8
           ,x"ffff" -- 73DA
           ,x"ffff" -- 73DC
           ,x"ffff" -- 73DE
           ,x"ffff" -- 73E0
           ,x"ffff" -- 73E2
           ,x"ffff" -- 73E4
           ,x"ffff" -- 73E6
           ,x"ffff" -- 73E8
           ,x"ffff" -- 73EA
           ,x"ffff" -- 73EC
           ,x"ffff" -- 73EE
           ,x"ffff" -- 73F0
           ,x"ffff" -- 73F2
           ,x"ffff" -- 73F4
           ,x"ffff" -- 73F6
           ,x"ffff" -- 73F8
           ,x"ffff" -- 73FA
           ,x"ffff" -- 73FC
           ,x"ffff" -- 73FE
           ,x"ffff" -- 7400
           ,x"ffff" -- 7402
           ,x"ffff" -- 7404
           ,x"ffff" -- 7406
           ,x"ffff" -- 7408
           ,x"ffff" -- 740A
           ,x"ffff" -- 740C
           ,x"ffff" -- 740E
           ,x"ffff" -- 7410
           ,x"ffff" -- 7412
           ,x"ffff" -- 7414
           ,x"ffff" -- 7416
           ,x"ffff" -- 7418
           ,x"ffff" -- 741A
           ,x"ffff" -- 741C
           ,x"ffff" -- 741E
           ,x"ffff" -- 7420
           ,x"ffff" -- 7422
           ,x"ffff" -- 7424
           ,x"ffff" -- 7426
           ,x"ffff" -- 7428
           ,x"ffff" -- 742A
           ,x"ffff" -- 742C
           ,x"ffff" -- 742E
           ,x"ffff" -- 7430
           ,x"ffff" -- 7432
           ,x"ffff" -- 7434
           ,x"ffff" -- 7436
           ,x"ffff" -- 7438
           ,x"ffff" -- 743A
           ,x"ffff" -- 743C
           ,x"ffff" -- 743E
           ,x"ffff" -- 7440
           ,x"ffff" -- 7442
           ,x"ffff" -- 7444
           ,x"ffff" -- 7446
           ,x"ffff" -- 7448
           ,x"ffff" -- 744A
           ,x"ffff" -- 744C
           ,x"ffff" -- 744E
           ,x"ffff" -- 7450
           ,x"ffff" -- 7452
           ,x"ffff" -- 7454
           ,x"ffff" -- 7456
           ,x"ffff" -- 7458
           ,x"ffff" -- 745A
           ,x"ffff" -- 745C
           ,x"ffff" -- 745E
           ,x"ffff" -- 7460
           ,x"ffff" -- 7462
           ,x"ffff" -- 7464
           ,x"ffff" -- 7466
           ,x"ffff" -- 7468
           ,x"ffff" -- 746A
           ,x"ffff" -- 746C
           ,x"ffff" -- 746E
           ,x"ffff" -- 7470
           ,x"ffff" -- 7472
           ,x"ffff" -- 7474
           ,x"ffff" -- 7476
           ,x"ffff" -- 7478
           ,x"ffff" -- 747A
           ,x"ffff" -- 747C
           ,x"ffff" -- 747E
           ,x"ffff" -- 7480
           ,x"ffff" -- 7482
           ,x"ffff" -- 7484
           ,x"ffff" -- 7486
           ,x"ffff" -- 7488
           ,x"ffff" -- 748A
           ,x"ffff" -- 748C
           ,x"ffff" -- 748E
           ,x"ffff" -- 7490
           ,x"ffff" -- 7492
           ,x"ffff" -- 7494
           ,x"ffff" -- 7496
           ,x"ffff" -- 7498
           ,x"ffff" -- 749A
           ,x"ffff" -- 749C
           ,x"ffff" -- 749E
           ,x"ffff" -- 74A0
           ,x"ffff" -- 74A2
           ,x"ffff" -- 74A4
           ,x"ffff" -- 74A6
           ,x"ffff" -- 74A8
           ,x"ffff" -- 74AA
           ,x"ffff" -- 74AC
           ,x"ffff" -- 74AE
           ,x"ffff" -- 74B0
           ,x"ffff" -- 74B2
           ,x"ffff" -- 74B4
           ,x"ffff" -- 74B6
           ,x"ffff" -- 74B8
           ,x"ffff" -- 74BA
           ,x"ffff" -- 74BC
           ,x"ffff" -- 74BE
           ,x"ffff" -- 74C0
           ,x"ffff" -- 74C2
           ,x"ffff" -- 74C4
           ,x"ffff" -- 74C6
           ,x"ffff" -- 74C8
           ,x"ffff" -- 74CA
           ,x"ffff" -- 74CC
           ,x"ffff" -- 74CE
           ,x"ffff" -- 74D0
           ,x"ffff" -- 74D2
           ,x"ffff" -- 74D4
           ,x"ffff" -- 74D6
           ,x"ffff" -- 74D8
           ,x"ffff" -- 74DA
           ,x"ffff" -- 74DC
           ,x"ffff" -- 74DE
           ,x"ffff" -- 74E0
           ,x"ffff" -- 74E2
           ,x"ffff" -- 74E4
           ,x"ffff" -- 74E6
           ,x"ffff" -- 74E8
           ,x"ffff" -- 74EA
           ,x"ffff" -- 74EC
           ,x"ffff" -- 74EE
           ,x"ffff" -- 74F0
           ,x"ffff" -- 74F2
           ,x"ffff" -- 74F4
           ,x"ffff" -- 74F6
           ,x"ffff" -- 74F8
           ,x"ffff" -- 74FA
           ,x"ffff" -- 74FC
           ,x"ffff" -- 74FE
           ,x"ffff" -- 7500
           ,x"ffff" -- 7502
           ,x"ffff" -- 7504
           ,x"ffff" -- 7506
           ,x"ffff" -- 7508
           ,x"ffff" -- 750A
           ,x"ffff" -- 750C
           ,x"ffff" -- 750E
           ,x"ffff" -- 7510
           ,x"ffff" -- 7512
           ,x"ffff" -- 7514
           ,x"ffff" -- 7516
           ,x"ffff" -- 7518
           ,x"ffff" -- 751A
           ,x"ffff" -- 751C
           ,x"ffff" -- 751E
           ,x"ffff" -- 7520
           ,x"ffff" -- 7522
           ,x"ffff" -- 7524
           ,x"ffff" -- 7526
           ,x"ffff" -- 7528
           ,x"ffff" -- 752A
           ,x"ffff" -- 752C
           ,x"ffff" -- 752E
           ,x"ffff" -- 7530
           ,x"ffff" -- 7532
           ,x"ffff" -- 7534
           ,x"ffff" -- 7536
           ,x"ffff" -- 7538
           ,x"ffff" -- 753A
           ,x"ffff" -- 753C
           ,x"ffff" -- 753E
           ,x"ffff" -- 7540
           ,x"ffff" -- 7542
           ,x"ffff" -- 7544
           ,x"ffff" -- 7546
           ,x"ffff" -- 7548
           ,x"ffff" -- 754A
           ,x"ffff" -- 754C
           ,x"ffff" -- 754E
           ,x"ffff" -- 7550
           ,x"ffff" -- 7552
           ,x"ffff" -- 7554
           ,x"ffff" -- 7556
           ,x"ffff" -- 7558
           ,x"ffff" -- 755A
           ,x"ffff" -- 755C
           ,x"ffff" -- 755E
           ,x"ffff" -- 7560
           ,x"ffff" -- 7562
           ,x"ffff" -- 7564
           ,x"ffff" -- 7566
           ,x"ffff" -- 7568
           ,x"ffff" -- 756A
           ,x"ffff" -- 756C
           ,x"ffff" -- 756E
           ,x"ffff" -- 7570
           ,x"ffff" -- 7572
           ,x"ffff" -- 7574
           ,x"ffff" -- 7576
           ,x"ffff" -- 7578
           ,x"ffff" -- 757A
           ,x"ffff" -- 757C
           ,x"ffff" -- 757E
           ,x"ffff" -- 7580
           ,x"ffff" -- 7582
           ,x"ffff" -- 7584
           ,x"ffff" -- 7586
           ,x"ffff" -- 7588
           ,x"ffff" -- 758A
           ,x"ffff" -- 758C
           ,x"ffff" -- 758E
           ,x"ffff" -- 7590
           ,x"ffff" -- 7592
           ,x"ffff" -- 7594
           ,x"ffff" -- 7596
           ,x"ffff" -- 7598
           ,x"ffff" -- 759A
           ,x"ffff" -- 759C
           ,x"ffff" -- 759E
           ,x"ffff" -- 75A0
           ,x"ffff" -- 75A2
           ,x"ffff" -- 75A4
           ,x"ffff" -- 75A6
           ,x"ffff" -- 75A8
           ,x"ffff" -- 75AA
           ,x"ffff" -- 75AC
           ,x"ffff" -- 75AE
           ,x"ffff" -- 75B0
           ,x"ffff" -- 75B2
           ,x"ffff" -- 75B4
           ,x"ffff" -- 75B6
           ,x"ffff" -- 75B8
           ,x"ffff" -- 75BA
           ,x"ffff" -- 75BC
           ,x"ffff" -- 75BE
           ,x"ffff" -- 75C0
           ,x"ffff" -- 75C2
           ,x"ffff" -- 75C4
           ,x"ffff" -- 75C6
           ,x"ffff" -- 75C8
           ,x"ffff" -- 75CA
           ,x"ffff" -- 75CC
           ,x"ffff" -- 75CE
           ,x"ffff" -- 75D0
           ,x"ffff" -- 75D2
           ,x"ffff" -- 75D4
           ,x"ffff" -- 75D6
           ,x"ffff" -- 75D8
           ,x"ffff" -- 75DA
           ,x"ffff" -- 75DC
           ,x"ffff" -- 75DE
           ,x"ffff" -- 75E0
           ,x"ffff" -- 75E2
           ,x"ffff" -- 75E4
           ,x"ffff" -- 75E6
           ,x"ffff" -- 75E8
           ,x"ffff" -- 75EA
           ,x"ffff" -- 75EC
           ,x"ffff" -- 75EE
           ,x"ffff" -- 75F0
           ,x"ffff" -- 75F2
           ,x"ffff" -- 75F4
           ,x"ffff" -- 75F6
           ,x"ffff" -- 75F8
           ,x"ffff" -- 75FA
           ,x"ffff" -- 75FC
           ,x"ffff" -- 75FE
           ,x"ffff" -- 7600
           ,x"ffff" -- 7602
           ,x"ffff" -- 7604
           ,x"ffff" -- 7606
           ,x"ffff" -- 7608
           ,x"ffff" -- 760A
           ,x"ffff" -- 760C
           ,x"ffff" -- 760E
           ,x"ffff" -- 7610
           ,x"ffff" -- 7612
           ,x"ffff" -- 7614
           ,x"ffff" -- 7616
           ,x"ffff" -- 7618
           ,x"ffff" -- 761A
           ,x"ffff" -- 761C
           ,x"ffff" -- 761E
           ,x"ffff" -- 7620
           ,x"ffff" -- 7622
           ,x"ffff" -- 7624
           ,x"ffff" -- 7626
           ,x"ffff" -- 7628
           ,x"ffff" -- 762A
           ,x"ffff" -- 762C
           ,x"ffff" -- 762E
           ,x"ffff" -- 7630
           ,x"ffff" -- 7632
           ,x"ffff" -- 7634
           ,x"ffff" -- 7636
           ,x"ffff" -- 7638
           ,x"ffff" -- 763A
           ,x"ffff" -- 763C
           ,x"ffff" -- 763E
           ,x"ffff" -- 7640
           ,x"ffff" -- 7642
           ,x"ffff" -- 7644
           ,x"ffff" -- 7646
           ,x"ffff" -- 7648
           ,x"ffff" -- 764A
           ,x"ffff" -- 764C
           ,x"ffff" -- 764E
           ,x"ffff" -- 7650
           ,x"ffff" -- 7652
           ,x"ffff" -- 7654
           ,x"ffff" -- 7656
           ,x"ffff" -- 7658
           ,x"ffff" -- 765A
           ,x"ffff" -- 765C
           ,x"ffff" -- 765E
           ,x"ffff" -- 7660
           ,x"ffff" -- 7662
           ,x"ffff" -- 7664
           ,x"ffff" -- 7666
           ,x"ffff" -- 7668
           ,x"ffff" -- 766A
           ,x"ffff" -- 766C
           ,x"ffff" -- 766E
           ,x"ffff" -- 7670
           ,x"ffff" -- 7672
           ,x"ffff" -- 7674
           ,x"ffff" -- 7676
           ,x"ffff" -- 7678
           ,x"ffff" -- 767A
           ,x"ffff" -- 767C
           ,x"ffff" -- 767E
           ,x"ffff" -- 7680
           ,x"ffff" -- 7682
           ,x"ffff" -- 7684
           ,x"ffff" -- 7686
           ,x"ffff" -- 7688
           ,x"ffff" -- 768A
           ,x"ffff" -- 768C
           ,x"ffff" -- 768E
           ,x"ffff" -- 7690
           ,x"ffff" -- 7692
           ,x"ffff" -- 7694
           ,x"ffff" -- 7696
           ,x"ffff" -- 7698
           ,x"ffff" -- 769A
           ,x"ffff" -- 769C
           ,x"ffff" -- 769E
           ,x"ffff" -- 76A0
           ,x"ffff" -- 76A2
           ,x"ffff" -- 76A4
           ,x"ffff" -- 76A6
           ,x"ffff" -- 76A8
           ,x"ffff" -- 76AA
           ,x"ffff" -- 76AC
           ,x"ffff" -- 76AE
           ,x"ffff" -- 76B0
           ,x"ffff" -- 76B2
           ,x"ffff" -- 76B4
           ,x"ffff" -- 76B6
           ,x"ffff" -- 76B8
           ,x"ffff" -- 76BA
           ,x"ffff" -- 76BC
           ,x"ffff" -- 76BE
           ,x"ffff" -- 76C0
           ,x"ffff" -- 76C2
           ,x"ffff" -- 76C4
           ,x"ffff" -- 76C6
           ,x"ffff" -- 76C8
           ,x"ffff" -- 76CA
           ,x"ffff" -- 76CC
           ,x"ffff" -- 76CE
           ,x"ffff" -- 76D0
           ,x"ffff" -- 76D2
           ,x"ffff" -- 76D4
           ,x"ffff" -- 76D6
           ,x"ffff" -- 76D8
           ,x"ffff" -- 76DA
           ,x"ffff" -- 76DC
           ,x"ffff" -- 76DE
           ,x"ffff" -- 76E0
           ,x"ffff" -- 76E2
           ,x"ffff" -- 76E4
           ,x"ffff" -- 76E6
           ,x"ffff" -- 76E8
           ,x"ffff" -- 76EA
           ,x"ffff" -- 76EC
           ,x"ffff" -- 76EE
           ,x"ffff" -- 76F0
           ,x"ffff" -- 76F2
           ,x"ffff" -- 76F4
           ,x"ffff" -- 76F6
           ,x"ffff" -- 76F8
           ,x"ffff" -- 76FA
           ,x"ffff" -- 76FC
           ,x"ffff" -- 76FE
           ,x"ffff" -- 7700
           ,x"ffff" -- 7702
           ,x"ffff" -- 7704
           ,x"ffff" -- 7706
           ,x"ffff" -- 7708
           ,x"ffff" -- 770A
           ,x"ffff" -- 770C
           ,x"ffff" -- 770E
           ,x"ffff" -- 7710
           ,x"ffff" -- 7712
           ,x"ffff" -- 7714
           ,x"ffff" -- 7716
           ,x"ffff" -- 7718
           ,x"ffff" -- 771A
           ,x"ffff" -- 771C
           ,x"ffff" -- 771E
           ,x"ffff" -- 7720
           ,x"ffff" -- 7722
           ,x"ffff" -- 7724
           ,x"ffff" -- 7726
           ,x"ffff" -- 7728
           ,x"ffff" -- 772A
           ,x"ffff" -- 772C
           ,x"ffff" -- 772E
           ,x"ffff" -- 7730
           ,x"ffff" -- 7732
           ,x"ffff" -- 7734
           ,x"ffff" -- 7736
           ,x"ffff" -- 7738
           ,x"ffff" -- 773A
           ,x"ffff" -- 773C
           ,x"ffff" -- 773E
           ,x"ffff" -- 7740
           ,x"ffff" -- 7742
           ,x"ffff" -- 7744
           ,x"ffff" -- 7746
           ,x"ffff" -- 7748
           ,x"ffff" -- 774A
           ,x"ffff" -- 774C
           ,x"ffff" -- 774E
           ,x"ffff" -- 7750
           ,x"ffff" -- 7752
           ,x"ffff" -- 7754
           ,x"ffff" -- 7756
           ,x"ffff" -- 7758
           ,x"ffff" -- 775A
           ,x"ffff" -- 775C
           ,x"ffff" -- 775E
           ,x"ffff" -- 7760
           ,x"ffff" -- 7762
           ,x"ffff" -- 7764
           ,x"ffff" -- 7766
           ,x"ffff" -- 7768
           ,x"ffff" -- 776A
           ,x"ffff" -- 776C
           ,x"ffff" -- 776E
           ,x"ffff" -- 7770
           ,x"ffff" -- 7772
           ,x"ffff" -- 7774
           ,x"ffff" -- 7776
           ,x"ffff" -- 7778
           ,x"ffff" -- 777A
           ,x"ffff" -- 777C
           ,x"ffff" -- 777E
           ,x"ffff" -- 7780
           ,x"ffff" -- 7782
           ,x"ffff" -- 7784
           ,x"ffff" -- 7786
           ,x"ffff" -- 7788
           ,x"ffff" -- 778A
           ,x"ffff" -- 778C
           ,x"ffff" -- 778E
           ,x"ffff" -- 7790
           ,x"ffff" -- 7792
           ,x"ffff" -- 7794
           ,x"ffff" -- 7796
           ,x"ffff" -- 7798
           ,x"ffff" -- 779A
           ,x"ffff" -- 779C
           ,x"ffff" -- 779E
           ,x"ffff" -- 77A0
           ,x"ffff" -- 77A2
           ,x"ffff" -- 77A4
           ,x"ffff" -- 77A6
           ,x"ffff" -- 77A8
           ,x"ffff" -- 77AA
           ,x"ffff" -- 77AC
           ,x"ffff" -- 77AE
           ,x"ffff" -- 77B0
           ,x"ffff" -- 77B2
           ,x"ffff" -- 77B4
           ,x"ffff" -- 77B6
           ,x"ffff" -- 77B8
           ,x"ffff" -- 77BA
           ,x"ffff" -- 77BC
           ,x"ffff" -- 77BE
           ,x"ffff" -- 77C0
           ,x"ffff" -- 77C2
           ,x"ffff" -- 77C4
           ,x"ffff" -- 77C6
           ,x"ffff" -- 77C8
           ,x"ffff" -- 77CA
           ,x"ffff" -- 77CC
           ,x"ffff" -- 77CE
           ,x"ffff" -- 77D0
           ,x"ffff" -- 77D2
           ,x"ffff" -- 77D4
           ,x"ffff" -- 77D6
           ,x"ffff" -- 77D8
           ,x"ffff" -- 77DA
           ,x"ffff" -- 77DC
           ,x"ffff" -- 77DE
           ,x"ffff" -- 77E0
           ,x"ffff" -- 77E2
           ,x"ffff" -- 77E4
           ,x"ffff" -- 77E6
           ,x"ffff" -- 77E8
           ,x"ffff" -- 77EA
           ,x"ffff" -- 77EC
           ,x"ffff" -- 77EE
           ,x"ffff" -- 77F0
           ,x"ffff" -- 77F2
           ,x"ffff" -- 77F4
           ,x"ffff" -- 77F6
           ,x"ffff" -- 77F8
           ,x"ffff" -- 77FA
           ,x"ffff" -- 77FC
           ,x"ffff" -- 77FE
           ,x"ffff" -- 7800
           ,x"ffff" -- 7802
           ,x"ffff" -- 7804
           ,x"ffff" -- 7806
           ,x"ffff" -- 7808
           ,x"ffff" -- 780A
           ,x"ffff" -- 780C
           ,x"ffff" -- 780E
           ,x"ffff" -- 7810
           ,x"ffff" -- 7812
           ,x"ffff" -- 7814
           ,x"ffff" -- 7816
           ,x"ffff" -- 7818
           ,x"ffff" -- 781A
           ,x"ffff" -- 781C
           ,x"ffff" -- 781E
           ,x"ffff" -- 7820
           ,x"ffff" -- 7822
           ,x"ffff" -- 7824
           ,x"ffff" -- 7826
           ,x"ffff" -- 7828
           ,x"ffff" -- 782A
           ,x"ffff" -- 782C
           ,x"ffff" -- 782E
           ,x"ffff" -- 7830
           ,x"ffff" -- 7832
           ,x"ffff" -- 7834
           ,x"ffff" -- 7836
           ,x"ffff" -- 7838
           ,x"ffff" -- 783A
           ,x"ffff" -- 783C
           ,x"ffff" -- 783E
           ,x"ffff" -- 7840
           ,x"ffff" -- 7842
           ,x"ffff" -- 7844
           ,x"ffff" -- 7846
           ,x"ffff" -- 7848
           ,x"ffff" -- 784A
           ,x"ffff" -- 784C
           ,x"ffff" -- 784E
           ,x"ffff" -- 7850
           ,x"ffff" -- 7852
           ,x"ffff" -- 7854
           ,x"ffff" -- 7856
           ,x"ffff" -- 7858
           ,x"ffff" -- 785A
           ,x"ffff" -- 785C
           ,x"ffff" -- 785E
           ,x"ffff" -- 7860
           ,x"ffff" -- 7862
           ,x"ffff" -- 7864
           ,x"ffff" -- 7866
           ,x"ffff" -- 7868
           ,x"ffff" -- 786A
           ,x"ffff" -- 786C
           ,x"ffff" -- 786E
           ,x"ffff" -- 7870
           ,x"ffff" -- 7872
           ,x"ffff" -- 7874
           ,x"ffff" -- 7876
           ,x"ffff" -- 7878
           ,x"ffff" -- 787A
           ,x"ffff" -- 787C
           ,x"ffff" -- 787E
           ,x"ffff" -- 7880
           ,x"ffff" -- 7882
           ,x"ffff" -- 7884
           ,x"ffff" -- 7886
           ,x"ffff" -- 7888
           ,x"ffff" -- 788A
           ,x"ffff" -- 788C
           ,x"ffff" -- 788E
           ,x"ffff" -- 7890
           ,x"ffff" -- 7892
           ,x"ffff" -- 7894
           ,x"ffff" -- 7896
           ,x"ffff" -- 7898
           ,x"ffff" -- 789A
           ,x"ffff" -- 789C
           ,x"ffff" -- 789E
           ,x"ffff" -- 78A0
           ,x"ffff" -- 78A2
           ,x"ffff" -- 78A4
           ,x"ffff" -- 78A6
           ,x"ffff" -- 78A8
           ,x"ffff" -- 78AA
           ,x"ffff" -- 78AC
           ,x"ffff" -- 78AE
           ,x"ffff" -- 78B0
           ,x"ffff" -- 78B2
           ,x"ffff" -- 78B4
           ,x"ffff" -- 78B6
           ,x"ffff" -- 78B8
           ,x"ffff" -- 78BA
           ,x"ffff" -- 78BC
           ,x"ffff" -- 78BE
           ,x"ffff" -- 78C0
           ,x"ffff" -- 78C2
           ,x"ffff" -- 78C4
           ,x"ffff" -- 78C6
           ,x"ffff" -- 78C8
           ,x"ffff" -- 78CA
           ,x"ffff" -- 78CC
           ,x"ffff" -- 78CE
           ,x"ffff" -- 78D0
           ,x"ffff" -- 78D2
           ,x"ffff" -- 78D4
           ,x"ffff" -- 78D6
           ,x"ffff" -- 78D8
           ,x"ffff" -- 78DA
           ,x"ffff" -- 78DC
           ,x"ffff" -- 78DE
           ,x"ffff" -- 78E0
           ,x"ffff" -- 78E2
           ,x"ffff" -- 78E4
           ,x"ffff" -- 78E6
           ,x"ffff" -- 78E8
           ,x"ffff" -- 78EA
           ,x"ffff" -- 78EC
           ,x"ffff" -- 78EE
           ,x"ffff" -- 78F0
           ,x"ffff" -- 78F2
           ,x"ffff" -- 78F4
           ,x"ffff" -- 78F6
           ,x"ffff" -- 78F8
           ,x"ffff" -- 78FA
           ,x"ffff" -- 78FC
           ,x"ffff" -- 78FE
           ,x"ffff" -- 7900
           ,x"ffff" -- 7902
           ,x"ffff" -- 7904
           ,x"ffff" -- 7906
           ,x"ffff" -- 7908
           ,x"ffff" -- 790A
           ,x"ffff" -- 790C
           ,x"ffff" -- 790E
           ,x"ffff" -- 7910
           ,x"ffff" -- 7912
           ,x"ffff" -- 7914
           ,x"ffff" -- 7916
           ,x"ffff" -- 7918
           ,x"ffff" -- 791A
           ,x"ffff" -- 791C
           ,x"ffff" -- 791E
           ,x"ffff" -- 7920
           ,x"ffff" -- 7922
           ,x"ffff" -- 7924
           ,x"ffff" -- 7926
           ,x"ffff" -- 7928
           ,x"ffff" -- 792A
           ,x"ffff" -- 792C
           ,x"ffff" -- 792E
           ,x"ffff" -- 7930
           ,x"ffff" -- 7932
           ,x"ffff" -- 7934
           ,x"ffff" -- 7936
           ,x"ffff" -- 7938
           ,x"ffff" -- 793A
           ,x"ffff" -- 793C
           ,x"ffff" -- 793E
           ,x"ffff" -- 7940
           ,x"ffff" -- 7942
           ,x"ffff" -- 7944
           ,x"ffff" -- 7946
           ,x"ffff" -- 7948
           ,x"ffff" -- 794A
           ,x"ffff" -- 794C
           ,x"ffff" -- 794E
           ,x"ffff" -- 7950
           ,x"ffff" -- 7952
           ,x"ffff" -- 7954
           ,x"ffff" -- 7956
           ,x"ffff" -- 7958
           ,x"ffff" -- 795A
           ,x"ffff" -- 795C
           ,x"ffff" -- 795E
           ,x"ffff" -- 7960
           ,x"ffff" -- 7962
           ,x"ffff" -- 7964
           ,x"ffff" -- 7966
           ,x"ffff" -- 7968
           ,x"ffff" -- 796A
           ,x"ffff" -- 796C
           ,x"ffff" -- 796E
           ,x"ffff" -- 7970
           ,x"ffff" -- 7972
           ,x"ffff" -- 7974
           ,x"ffff" -- 7976
           ,x"ffff" -- 7978
           ,x"ffff" -- 797A
           ,x"ffff" -- 797C
           ,x"ffff" -- 797E
           ,x"ffff" -- 7980
           ,x"ffff" -- 7982
           ,x"ffff" -- 7984
           ,x"ffff" -- 7986
           ,x"ffff" -- 7988
           ,x"ffff" -- 798A
           ,x"ffff" -- 798C
           ,x"ffff" -- 798E
           ,x"ffff" -- 7990
           ,x"ffff" -- 7992
           ,x"ffff" -- 7994
           ,x"ffff" -- 7996
           ,x"ffff" -- 7998
           ,x"ffff" -- 799A
           ,x"ffff" -- 799C
           ,x"ffff" -- 799E
           ,x"ffff" -- 79A0
           ,x"ffff" -- 79A2
           ,x"ffff" -- 79A4
           ,x"ffff" -- 79A6
           ,x"ffff" -- 79A8
           ,x"ffff" -- 79AA
           ,x"ffff" -- 79AC
           ,x"ffff" -- 79AE
           ,x"ffff" -- 79B0
           ,x"ffff" -- 79B2
           ,x"ffff" -- 79B4
           ,x"ffff" -- 79B6
           ,x"ffff" -- 79B8
           ,x"ffff" -- 79BA
           ,x"ffff" -- 79BC
           ,x"ffff" -- 79BE
           ,x"ffff" -- 79C0
           ,x"ffff" -- 79C2
           ,x"ffff" -- 79C4
           ,x"ffff" -- 79C6
           ,x"ffff" -- 79C8
           ,x"ffff" -- 79CA
           ,x"ffff" -- 79CC
           ,x"ffff" -- 79CE
           ,x"ffff" -- 79D0
           ,x"ffff" -- 79D2
           ,x"ffff" -- 79D4
           ,x"ffff" -- 79D6
           ,x"ffff" -- 79D8
           ,x"ffff" -- 79DA
           ,x"ffff" -- 79DC
           ,x"ffff" -- 79DE
           ,x"ffff" -- 79E0
           ,x"ffff" -- 79E2
           ,x"ffff" -- 79E4
           ,x"ffff" -- 79E6
           ,x"ffff" -- 79E8
           ,x"ffff" -- 79EA
           ,x"ffff" -- 79EC
           ,x"ffff" -- 79EE
           ,x"ffff" -- 79F0
           ,x"ffff" -- 79F2
           ,x"ffff" -- 79F4
           ,x"ffff" -- 79F6
           ,x"ffff" -- 79F8
           ,x"ffff" -- 79FA
           ,x"ffff" -- 79FC
           ,x"ffff" -- 79FE
           ,x"ffff" -- 7A00
           ,x"ffff" -- 7A02
           ,x"ffff" -- 7A04
           ,x"ffff" -- 7A06
           ,x"ffff" -- 7A08
           ,x"ffff" -- 7A0A
           ,x"ffff" -- 7A0C
           ,x"ffff" -- 7A0E
           ,x"ffff" -- 7A10
           ,x"ffff" -- 7A12
           ,x"ffff" -- 7A14
           ,x"ffff" -- 7A16
           ,x"ffff" -- 7A18
           ,x"ffff" -- 7A1A
           ,x"ffff" -- 7A1C
           ,x"ffff" -- 7A1E
           ,x"ffff" -- 7A20
           ,x"ffff" -- 7A22
           ,x"ffff" -- 7A24
           ,x"ffff" -- 7A26
           ,x"ffff" -- 7A28
           ,x"ffff" -- 7A2A
           ,x"ffff" -- 7A2C
           ,x"ffff" -- 7A2E
           ,x"ffff" -- 7A30
           ,x"ffff" -- 7A32
           ,x"ffff" -- 7A34
           ,x"ffff" -- 7A36
           ,x"ffff" -- 7A38
           ,x"ffff" -- 7A3A
           ,x"ffff" -- 7A3C
           ,x"ffff" -- 7A3E
           ,x"ffff" -- 7A40
           ,x"ffff" -- 7A42
           ,x"ffff" -- 7A44
           ,x"ffff" -- 7A46
           ,x"ffff" -- 7A48
           ,x"ffff" -- 7A4A
           ,x"ffff" -- 7A4C
           ,x"ffff" -- 7A4E
           ,x"ffff" -- 7A50
           ,x"ffff" -- 7A52
           ,x"ffff" -- 7A54
           ,x"ffff" -- 7A56
           ,x"ffff" -- 7A58
           ,x"ffff" -- 7A5A
           ,x"ffff" -- 7A5C
           ,x"ffff" -- 7A5E
           ,x"ffff" -- 7A60
           ,x"ffff" -- 7A62
           ,x"ffff" -- 7A64
           ,x"ffff" -- 7A66
           ,x"ffff" -- 7A68
           ,x"ffff" -- 7A6A
           ,x"ffff" -- 7A6C
           ,x"ffff" -- 7A6E
           ,x"ffff" -- 7A70
           ,x"ffff" -- 7A72
           ,x"ffff" -- 7A74
           ,x"ffff" -- 7A76
           ,x"ffff" -- 7A78
           ,x"ffff" -- 7A7A
           ,x"ffff" -- 7A7C
           ,x"ffff" -- 7A7E
           ,x"ffff" -- 7A80
           ,x"ffff" -- 7A82
           ,x"ffff" -- 7A84
           ,x"ffff" -- 7A86
           ,x"ffff" -- 7A88
           ,x"ffff" -- 7A8A
           ,x"ffff" -- 7A8C
           ,x"ffff" -- 7A8E
           ,x"ffff" -- 7A90
           ,x"ffff" -- 7A92
           ,x"ffff" -- 7A94
           ,x"ffff" -- 7A96
           ,x"ffff" -- 7A98
           ,x"ffff" -- 7A9A
           ,x"ffff" -- 7A9C
           ,x"ffff" -- 7A9E
           ,x"ffff" -- 7AA0
           ,x"ffff" -- 7AA2
           ,x"ffff" -- 7AA4
           ,x"ffff" -- 7AA6
           ,x"ffff" -- 7AA8
           ,x"ffff" -- 7AAA
           ,x"ffff" -- 7AAC
           ,x"ffff" -- 7AAE
           ,x"ffff" -- 7AB0
           ,x"ffff" -- 7AB2
           ,x"ffff" -- 7AB4
           ,x"ffff" -- 7AB6
           ,x"ffff" -- 7AB8
           ,x"ffff" -- 7ABA
           ,x"ffff" -- 7ABC
           ,x"ffff" -- 7ABE
           ,x"ffff" -- 7AC0
           ,x"ffff" -- 7AC2
           ,x"ffff" -- 7AC4
           ,x"ffff" -- 7AC6
           ,x"ffff" -- 7AC8
           ,x"ffff" -- 7ACA
           ,x"ffff" -- 7ACC
           ,x"ffff" -- 7ACE
           ,x"ffff" -- 7AD0
           ,x"ffff" -- 7AD2
           ,x"ffff" -- 7AD4
           ,x"ffff" -- 7AD6
           ,x"ffff" -- 7AD8
           ,x"ffff" -- 7ADA
           ,x"ffff" -- 7ADC
           ,x"ffff" -- 7ADE
           ,x"ffff" -- 7AE0
           ,x"ffff" -- 7AE2
           ,x"ffff" -- 7AE4
           ,x"ffff" -- 7AE6
           ,x"ffff" -- 7AE8
           ,x"ffff" -- 7AEA
           ,x"ffff" -- 7AEC
           ,x"ffff" -- 7AEE
           ,x"ffff" -- 7AF0
           ,x"ffff" -- 7AF2
           ,x"ffff" -- 7AF4
           ,x"ffff" -- 7AF6
           ,x"ffff" -- 7AF8
           ,x"ffff" -- 7AFA
           ,x"ffff" -- 7AFC
           ,x"ffff" -- 7AFE
           ,x"ffff" -- 7B00
           ,x"ffff" -- 7B02
           ,x"ffff" -- 7B04
           ,x"ffff" -- 7B06
           ,x"ffff" -- 7B08
           ,x"ffff" -- 7B0A
           ,x"ffff" -- 7B0C
           ,x"ffff" -- 7B0E
           ,x"ffff" -- 7B10
           ,x"ffff" -- 7B12
           ,x"ffff" -- 7B14
           ,x"ffff" -- 7B16
           ,x"ffff" -- 7B18
           ,x"ffff" -- 7B1A
           ,x"ffff" -- 7B1C
           ,x"ffff" -- 7B1E
           ,x"ffff" -- 7B20
           ,x"ffff" -- 7B22
           ,x"ffff" -- 7B24
           ,x"ffff" -- 7B26
           ,x"ffff" -- 7B28
           ,x"ffff" -- 7B2A
           ,x"ffff" -- 7B2C
           ,x"ffff" -- 7B2E
           ,x"ffff" -- 7B30
           ,x"ffff" -- 7B32
           ,x"ffff" -- 7B34
           ,x"ffff" -- 7B36
           ,x"ffff" -- 7B38
           ,x"ffff" -- 7B3A
           ,x"ffff" -- 7B3C
           ,x"ffff" -- 7B3E
           ,x"ffff" -- 7B40
           ,x"ffff" -- 7B42
           ,x"ffff" -- 7B44
           ,x"ffff" -- 7B46
           ,x"ffff" -- 7B48
           ,x"ffff" -- 7B4A
           ,x"ffff" -- 7B4C
           ,x"ffff" -- 7B4E
           ,x"ffff" -- 7B50
           ,x"ffff" -- 7B52
           ,x"ffff" -- 7B54
           ,x"ffff" -- 7B56
           ,x"ffff" -- 7B58
           ,x"ffff" -- 7B5A
           ,x"ffff" -- 7B5C
           ,x"ffff" -- 7B5E
           ,x"ffff" -- 7B60
           ,x"ffff" -- 7B62
           ,x"ffff" -- 7B64
           ,x"ffff" -- 7B66
           ,x"ffff" -- 7B68
           ,x"ffff" -- 7B6A
           ,x"ffff" -- 7B6C
           ,x"ffff" -- 7B6E
           ,x"ffff" -- 7B70
           ,x"ffff" -- 7B72
           ,x"ffff" -- 7B74
           ,x"ffff" -- 7B76
           ,x"ffff" -- 7B78
           ,x"ffff" -- 7B7A
           ,x"ffff" -- 7B7C
           ,x"ffff" -- 7B7E
           ,x"ffff" -- 7B80
           ,x"ffff" -- 7B82
           ,x"ffff" -- 7B84
           ,x"ffff" -- 7B86
           ,x"ffff" -- 7B88
           ,x"ffff" -- 7B8A
           ,x"ffff" -- 7B8C
           ,x"ffff" -- 7B8E
           ,x"ffff" -- 7B90
           ,x"ffff" -- 7B92
           ,x"ffff" -- 7B94
           ,x"ffff" -- 7B96
           ,x"ffff" -- 7B98
           ,x"ffff" -- 7B9A
           ,x"ffff" -- 7B9C
           ,x"ffff" -- 7B9E
           ,x"ffff" -- 7BA0
           ,x"ffff" -- 7BA2
           ,x"ffff" -- 7BA4
           ,x"ffff" -- 7BA6
           ,x"ffff" -- 7BA8
           ,x"ffff" -- 7BAA
           ,x"ffff" -- 7BAC
           ,x"ffff" -- 7BAE
           ,x"ffff" -- 7BB0
           ,x"ffff" -- 7BB2
           ,x"ffff" -- 7BB4
           ,x"ffff" -- 7BB6
           ,x"ffff" -- 7BB8
           ,x"ffff" -- 7BBA
           ,x"ffff" -- 7BBC
           ,x"ffff" -- 7BBE
           ,x"ffff" -- 7BC0
           ,x"ffff" -- 7BC2
           ,x"ffff" -- 7BC4
           ,x"ffff" -- 7BC6
           ,x"ffff" -- 7BC8
           ,x"ffff" -- 7BCA
           ,x"ffff" -- 7BCC
           ,x"ffff" -- 7BCE
           ,x"ffff" -- 7BD0
           ,x"ffff" -- 7BD2
           ,x"ffff" -- 7BD4
           ,x"ffff" -- 7BD6
           ,x"ffff" -- 7BD8
           ,x"ffff" -- 7BDA
           ,x"ffff" -- 7BDC
           ,x"ffff" -- 7BDE
           ,x"ffff" -- 7BE0
           ,x"ffff" -- 7BE2
           ,x"ffff" -- 7BE4
           ,x"ffff" -- 7BE6
           ,x"ffff" -- 7BE8
           ,x"ffff" -- 7BEA
           ,x"ffff" -- 7BEC
           ,x"ffff" -- 7BEE
           ,x"ffff" -- 7BF0
           ,x"ffff" -- 7BF2
           ,x"ffff" -- 7BF4
           ,x"ffff" -- 7BF6
           ,x"ffff" -- 7BF8
           ,x"ffff" -- 7BFA
           ,x"ffff" -- 7BFC
           ,x"ffff" -- 7BFE
           ,x"ffff" -- 7C00
           ,x"ffff" -- 7C02
           ,x"ffff" -- 7C04
           ,x"ffff" -- 7C06
           ,x"ffff" -- 7C08
           ,x"ffff" -- 7C0A
           ,x"ffff" -- 7C0C
           ,x"ffff" -- 7C0E
           ,x"ffff" -- 7C10
           ,x"ffff" -- 7C12
           ,x"ffff" -- 7C14
           ,x"ffff" -- 7C16
           ,x"ffff" -- 7C18
           ,x"ffff" -- 7C1A
           ,x"ffff" -- 7C1C
           ,x"ffff" -- 7C1E
           ,x"ffff" -- 7C20
           ,x"ffff" -- 7C22
           ,x"ffff" -- 7C24
           ,x"ffff" -- 7C26
           ,x"ffff" -- 7C28
           ,x"ffff" -- 7C2A
           ,x"ffff" -- 7C2C
           ,x"ffff" -- 7C2E
           ,x"ffff" -- 7C30
           ,x"ffff" -- 7C32
           ,x"ffff" -- 7C34
           ,x"ffff" -- 7C36
           ,x"ffff" -- 7C38
           ,x"ffff" -- 7C3A
           ,x"ffff" -- 7C3C
           ,x"ffff" -- 7C3E
           ,x"ffff" -- 7C40
           ,x"ffff" -- 7C42
           ,x"ffff" -- 7C44
           ,x"ffff" -- 7C46
           ,x"ffff" -- 7C48
           ,x"ffff" -- 7C4A
           ,x"ffff" -- 7C4C
           ,x"ffff" -- 7C4E
           ,x"ffff" -- 7C50
           ,x"ffff" -- 7C52
           ,x"ffff" -- 7C54
           ,x"ffff" -- 7C56
           ,x"ffff" -- 7C58
           ,x"ffff" -- 7C5A
           ,x"ffff" -- 7C5C
           ,x"ffff" -- 7C5E
           ,x"ffff" -- 7C60
           ,x"ffff" -- 7C62
           ,x"ffff" -- 7C64
           ,x"ffff" -- 7C66
           ,x"ffff" -- 7C68
           ,x"ffff" -- 7C6A
           ,x"ffff" -- 7C6C
           ,x"ffff" -- 7C6E
           ,x"ffff" -- 7C70
           ,x"ffff" -- 7C72
           ,x"ffff" -- 7C74
           ,x"ffff" -- 7C76
           ,x"ffff" -- 7C78
           ,x"ffff" -- 7C7A
           ,x"ffff" -- 7C7C
           ,x"ffff" -- 7C7E
           ,x"ffff" -- 7C80
           ,x"ffff" -- 7C82
           ,x"ffff" -- 7C84
           ,x"ffff" -- 7C86
           ,x"ffff" -- 7C88
           ,x"ffff" -- 7C8A
           ,x"ffff" -- 7C8C
           ,x"ffff" -- 7C8E
           ,x"ffff" -- 7C90
           ,x"ffff" -- 7C92
           ,x"ffff" -- 7C94
           ,x"ffff" -- 7C96
           ,x"ffff" -- 7C98
           ,x"ffff" -- 7C9A
           ,x"ffff" -- 7C9C
           ,x"ffff" -- 7C9E
           ,x"ffff" -- 7CA0
           ,x"ffff" -- 7CA2
           ,x"ffff" -- 7CA4
           ,x"ffff" -- 7CA6
           ,x"ffff" -- 7CA8
           ,x"ffff" -- 7CAA
           ,x"ffff" -- 7CAC
           ,x"ffff" -- 7CAE
           ,x"ffff" -- 7CB0
           ,x"ffff" -- 7CB2
           ,x"ffff" -- 7CB4
           ,x"ffff" -- 7CB6
           ,x"ffff" -- 7CB8
           ,x"ffff" -- 7CBA
           ,x"ffff" -- 7CBC
           ,x"ffff" -- 7CBE
           ,x"ffff" -- 7CC0
           ,x"ffff" -- 7CC2
           ,x"ffff" -- 7CC4
           ,x"ffff" -- 7CC6
           ,x"ffff" -- 7CC8
           ,x"ffff" -- 7CCA
           ,x"ffff" -- 7CCC
           ,x"ffff" -- 7CCE
           ,x"ffff" -- 7CD0
           ,x"ffff" -- 7CD2
           ,x"ffff" -- 7CD4
           ,x"ffff" -- 7CD6
           ,x"ffff" -- 7CD8
           ,x"ffff" -- 7CDA
           ,x"ffff" -- 7CDC
           ,x"ffff" -- 7CDE
           ,x"ffff" -- 7CE0
           ,x"ffff" -- 7CE2
           ,x"ffff" -- 7CE4
           ,x"ffff" -- 7CE6
           ,x"ffff" -- 7CE8
           ,x"ffff" -- 7CEA
           ,x"ffff" -- 7CEC
           ,x"ffff" -- 7CEE
           ,x"ffff" -- 7CF0
           ,x"ffff" -- 7CF2
           ,x"ffff" -- 7CF4
           ,x"ffff" -- 7CF6
           ,x"ffff" -- 7CF8
           ,x"ffff" -- 7CFA
           ,x"ffff" -- 7CFC
           ,x"ffff" -- 7CFE
           ,x"ffff" -- 7D00
           ,x"ffff" -- 7D02
           ,x"ffff" -- 7D04
           ,x"ffff" -- 7D06
           ,x"ffff" -- 7D08
           ,x"ffff" -- 7D0A
           ,x"ffff" -- 7D0C
           ,x"ffff" -- 7D0E
           ,x"ffff" -- 7D10
           ,x"ffff" -- 7D12
           ,x"ffff" -- 7D14
           ,x"ffff" -- 7D16
           ,x"ffff" -- 7D18
           ,x"ffff" -- 7D1A
           ,x"ffff" -- 7D1C
           ,x"ffff" -- 7D1E
           ,x"ffff" -- 7D20
           ,x"ffff" -- 7D22
           ,x"ffff" -- 7D24
           ,x"ffff" -- 7D26
           ,x"ffff" -- 7D28
           ,x"ffff" -- 7D2A
           ,x"ffff" -- 7D2C
           ,x"ffff" -- 7D2E
           ,x"ffff" -- 7D30
           ,x"ffff" -- 7D32
           ,x"ffff" -- 7D34
           ,x"ffff" -- 7D36
           ,x"ffff" -- 7D38
           ,x"ffff" -- 7D3A
           ,x"ffff" -- 7D3C
           ,x"ffff" -- 7D3E
           ,x"ffff" -- 7D40
           ,x"ffff" -- 7D42
           ,x"ffff" -- 7D44
           ,x"ffff" -- 7D46
           ,x"ffff" -- 7D48
           ,x"ffff" -- 7D4A
           ,x"ffff" -- 7D4C
           ,x"ffff" -- 7D4E
           ,x"ffff" -- 7D50
           ,x"ffff" -- 7D52
           ,x"ffff" -- 7D54
           ,x"ffff" -- 7D56
           ,x"ffff" -- 7D58
           ,x"ffff" -- 7D5A
           ,x"ffff" -- 7D5C
           ,x"ffff" -- 7D5E
           ,x"ffff" -- 7D60
           ,x"ffff" -- 7D62
           ,x"ffff" -- 7D64
           ,x"ffff" -- 7D66
           ,x"ffff" -- 7D68
           ,x"ffff" -- 7D6A
           ,x"ffff" -- 7D6C
           ,x"ffff" -- 7D6E
           ,x"ffff" -- 7D70
           ,x"ffff" -- 7D72
           ,x"ffff" -- 7D74
           ,x"ffff" -- 7D76
           ,x"ffff" -- 7D78
           ,x"ffff" -- 7D7A
           ,x"ffff" -- 7D7C
           ,x"ffff" -- 7D7E
           ,x"ffff" -- 7D80
           ,x"ffff" -- 7D82
           ,x"ffff" -- 7D84
           ,x"ffff" -- 7D86
           ,x"ffff" -- 7D88
           ,x"ffff" -- 7D8A
           ,x"ffff" -- 7D8C
           ,x"ffff" -- 7D8E
           ,x"ffff" -- 7D90
           ,x"ffff" -- 7D92
           ,x"ffff" -- 7D94
           ,x"ffff" -- 7D96
           ,x"ffff" -- 7D98
           ,x"ffff" -- 7D9A
           ,x"ffff" -- 7D9C
           ,x"ffff" -- 7D9E
           ,x"ffff" -- 7DA0
           ,x"ffff" -- 7DA2
           ,x"ffff" -- 7DA4
           ,x"ffff" -- 7DA6
           ,x"ffff" -- 7DA8
           ,x"ffff" -- 7DAA
           ,x"ffff" -- 7DAC
           ,x"ffff" -- 7DAE
           ,x"ffff" -- 7DB0
           ,x"ffff" -- 7DB2
           ,x"ffff" -- 7DB4
           ,x"ffff" -- 7DB6
           ,x"ffff" -- 7DB8
           ,x"ffff" -- 7DBA
           ,x"ffff" -- 7DBC
           ,x"ffff" -- 7DBE
           ,x"ffff" -- 7DC0
           ,x"ffff" -- 7DC2
           ,x"ffff" -- 7DC4
           ,x"ffff" -- 7DC6
           ,x"ffff" -- 7DC8
           ,x"ffff" -- 7DCA
           ,x"ffff" -- 7DCC
           ,x"ffff" -- 7DCE
           ,x"ffff" -- 7DD0
           ,x"ffff" -- 7DD2
           ,x"ffff" -- 7DD4
           ,x"ffff" -- 7DD6
           ,x"ffff" -- 7DD8
           ,x"ffff" -- 7DDA
           ,x"ffff" -- 7DDC
           ,x"ffff" -- 7DDE
           ,x"ffff" -- 7DE0
           ,x"ffff" -- 7DE2
           ,x"ffff" -- 7DE4
           ,x"ffff" -- 7DE6
           ,x"ffff" -- 7DE8
           ,x"ffff" -- 7DEA
           ,x"ffff" -- 7DEC
           ,x"ffff" -- 7DEE
           ,x"ffff" -- 7DF0
           ,x"ffff" -- 7DF2
           ,x"ffff" -- 7DF4
           ,x"ffff" -- 7DF6
           ,x"ffff" -- 7DF8
           ,x"ffff" -- 7DFA
           ,x"ffff" -- 7DFC
           ,x"ffff" -- 7DFE
           ,x"ffff" -- 7E00
           ,x"ffff" -- 7E02
           ,x"ffff" -- 7E04
           ,x"ffff" -- 7E06
           ,x"ffff" -- 7E08
           ,x"ffff" -- 7E0A
           ,x"ffff" -- 7E0C
           ,x"ffff" -- 7E0E
           ,x"ffff" -- 7E10
           ,x"ffff" -- 7E12
           ,x"ffff" -- 7E14
           ,x"ffff" -- 7E16
           ,x"ffff" -- 7E18
           ,x"ffff" -- 7E1A
           ,x"ffff" -- 7E1C
           ,x"ffff" -- 7E1E
           ,x"ffff" -- 7E20
           ,x"ffff" -- 7E22
           ,x"ffff" -- 7E24
           ,x"ffff" -- 7E26
           ,x"ffff" -- 7E28
           ,x"ffff" -- 7E2A
           ,x"ffff" -- 7E2C
           ,x"ffff" -- 7E2E
           ,x"ffff" -- 7E30
           ,x"ffff" -- 7E32
           ,x"ffff" -- 7E34
           ,x"ffff" -- 7E36
           ,x"ffff" -- 7E38
           ,x"ffff" -- 7E3A
           ,x"ffff" -- 7E3C
           ,x"ffff" -- 7E3E
           ,x"ffff" -- 7E40
           ,x"ffff" -- 7E42
           ,x"ffff" -- 7E44
           ,x"ffff" -- 7E46
           ,x"ffff" -- 7E48
           ,x"ffff" -- 7E4A
           ,x"ffff" -- 7E4C
           ,x"ffff" -- 7E4E
           ,x"ffff" -- 7E50
           ,x"ffff" -- 7E52
           ,x"ffff" -- 7E54
           ,x"ffff" -- 7E56
           ,x"ffff" -- 7E58
           ,x"ffff" -- 7E5A
           ,x"ffff" -- 7E5C
           ,x"ffff" -- 7E5E
           ,x"ffff" -- 7E60
           ,x"ffff" -- 7E62
           ,x"ffff" -- 7E64
           ,x"ffff" -- 7E66
           ,x"ffff" -- 7E68
           ,x"ffff" -- 7E6A
           ,x"ffff" -- 7E6C
           ,x"ffff" -- 7E6E
           ,x"ffff" -- 7E70
           ,x"ffff" -- 7E72
           ,x"ffff" -- 7E74
           ,x"ffff" -- 7E76
           ,x"ffff" -- 7E78
           ,x"ffff" -- 7E7A
           ,x"ffff" -- 7E7C
           ,x"ffff" -- 7E7E
           ,x"ffff" -- 7E80
           ,x"ffff" -- 7E82
           ,x"ffff" -- 7E84
           ,x"ffff" -- 7E86
           ,x"ffff" -- 7E88
           ,x"ffff" -- 7E8A
           ,x"ffff" -- 7E8C
           ,x"ffff" -- 7E8E
           ,x"ffff" -- 7E90
           ,x"ffff" -- 7E92
           ,x"ffff" -- 7E94
           ,x"ffff" -- 7E96
           ,x"ffff" -- 7E98
           ,x"ffff" -- 7E9A
           ,x"ffff" -- 7E9C
           ,x"ffff" -- 7E9E
           ,x"ffff" -- 7EA0
           ,x"ffff" -- 7EA2
           ,x"ffff" -- 7EA4
           ,x"ffff" -- 7EA6
           ,x"ffff" -- 7EA8
           ,x"ffff" -- 7EAA
           ,x"ffff" -- 7EAC
           ,x"ffff" -- 7EAE
           ,x"ffff" -- 7EB0
           ,x"ffff" -- 7EB2
           ,x"ffff" -- 7EB4
           ,x"ffff" -- 7EB6
           ,x"ffff" -- 7EB8
           ,x"ffff" -- 7EBA
           ,x"ffff" -- 7EBC
           ,x"ffff" -- 7EBE
           ,x"ffff" -- 7EC0
           ,x"ffff" -- 7EC2
           ,x"ffff" -- 7EC4
           ,x"ffff" -- 7EC6
           ,x"ffff" -- 7EC8
           ,x"ffff" -- 7ECA
           ,x"ffff" -- 7ECC
           ,x"ffff" -- 7ECE
           ,x"ffff" -- 7ED0
           ,x"ffff" -- 7ED2
           ,x"ffff" -- 7ED4
           ,x"ffff" -- 7ED6
           ,x"ffff" -- 7ED8
           ,x"ffff" -- 7EDA
           ,x"ffff" -- 7EDC
           ,x"ffff" -- 7EDE
           ,x"ffff" -- 7EE0
           ,x"ffff" -- 7EE2
           ,x"ffff" -- 7EE4
           ,x"ffff" -- 7EE6
           ,x"ffff" -- 7EE8
           ,x"ffff" -- 7EEA
           ,x"ffff" -- 7EEC
           ,x"ffff" -- 7EEE
           ,x"ffff" -- 7EF0
           ,x"ffff" -- 7EF2
           ,x"ffff" -- 7EF4
           ,x"ffff" -- 7EF6
           ,x"ffff" -- 7EF8
           ,x"ffff" -- 7EFA
           ,x"ffff" -- 7EFC
           ,x"ffff" -- 7EFE
           ,x"ffff" -- 7F00
           ,x"ffff" -- 7F02
           ,x"ffff" -- 7F04
           ,x"ffff" -- 7F06
           ,x"ffff" -- 7F08
           ,x"ffff" -- 7F0A
           ,x"ffff" -- 7F0C
           ,x"ffff" -- 7F0E
           ,x"ffff" -- 7F10
           ,x"ffff" -- 7F12
           ,x"ffff" -- 7F14
           ,x"ffff" -- 7F16
           ,x"ffff" -- 7F18
           ,x"ffff" -- 7F1A
           ,x"ffff" -- 7F1C
           ,x"ffff" -- 7F1E
           ,x"ffff" -- 7F20
           ,x"ffff" -- 7F22
           ,x"ffff" -- 7F24
           ,x"ffff" -- 7F26
           ,x"ffff" -- 7F28
           ,x"ffff" -- 7F2A
           ,x"ffff" -- 7F2C
           ,x"ffff" -- 7F2E
           ,x"ffff" -- 7F30
           ,x"ffff" -- 7F32
           ,x"ffff" -- 7F34
           ,x"ffff" -- 7F36
           ,x"ffff" -- 7F38
           ,x"ffff" -- 7F3A
           ,x"ffff" -- 7F3C
           ,x"ffff" -- 7F3E
           ,x"ffff" -- 7F40
           ,x"ffff" -- 7F42
           ,x"ffff" -- 7F44
           ,x"ffff" -- 7F46
           ,x"ffff" -- 7F48
           ,x"ffff" -- 7F4A
           ,x"ffff" -- 7F4C
           ,x"ffff" -- 7F4E
           ,x"ffff" -- 7F50
           ,x"ffff" -- 7F52
           ,x"ffff" -- 7F54
           ,x"ffff" -- 7F56
           ,x"ffff" -- 7F58
           ,x"ffff" -- 7F5A
           ,x"ffff" -- 7F5C
           ,x"ffff" -- 7F5E
           ,x"ffff" -- 7F60
           ,x"ffff" -- 7F62
           ,x"ffff" -- 7F64
           ,x"ffff" -- 7F66
           ,x"ffff" -- 7F68
           ,x"ffff" -- 7F6A
           ,x"ffff" -- 7F6C
           ,x"ffff" -- 7F6E
           ,x"ffff" -- 7F70
           ,x"ffff" -- 7F72
           ,x"ffff" -- 7F74
           ,x"ffff" -- 7F76
           ,x"ffff" -- 7F78
           ,x"ffff" -- 7F7A
           ,x"ffff" -- 7F7C
           ,x"ffff" -- 7F7E
           ,x"ffff" -- 7F80
           ,x"ffff" -- 7F82
           ,x"ffff" -- 7F84
           ,x"ffff" -- 7F86
           ,x"ffff" -- 7F88
           ,x"ffff" -- 7F8A
           ,x"ffff" -- 7F8C
           ,x"ffff" -- 7F8E
           ,x"ffff" -- 7F90
           ,x"ffff" -- 7F92
           ,x"ffff" -- 7F94
           ,x"ffff" -- 7F96
           ,x"ffff" -- 7F98
           ,x"ffff" -- 7F9A
           ,x"ffff" -- 7F9C
           ,x"ffff" -- 7F9E
           ,x"ffff" -- 7FA0
           ,x"ffff" -- 7FA2
           ,x"ffff" -- 7FA4
           ,x"ffff" -- 7FA6
           ,x"ffff" -- 7FA8
           ,x"ffff" -- 7FAA
           ,x"ffff" -- 7FAC
           ,x"ffff" -- 7FAE
           ,x"ffff" -- 7FB0
           ,x"ffff" -- 7FB2
           ,x"ffff" -- 7FB4
           ,x"ffff" -- 7FB6
           ,x"ffff" -- 7FB8
           ,x"ffff" -- 7FBA
           ,x"ffff" -- 7FBC
           ,x"ffff" -- 7FBE
           ,x"ffff" -- 7FC0
           ,x"ffff" -- 7FC2
           ,x"ffff" -- 7FC4
           ,x"ffff" -- 7FC6
           ,x"ffff" -- 7FC8
           ,x"ffff" -- 7FCA
           ,x"ffff" -- 7FCC
           ,x"ffff" -- 7FCE
           ,x"ffff" -- 7FD0
           ,x"ffff" -- 7FD2
           ,x"ffff" -- 7FD4
           ,x"ffff" -- 7FD6
           ,x"ffff" -- 7FD8
           ,x"ffff" -- 7FDA
           ,x"ffff" -- 7FDC
           ,x"ffff" -- 7FDE
           ,x"ffff" -- 7FE0
           ,x"ffff" -- 7FE2
           ,x"ffff" -- 7FE4
           ,x"ffff" -- 7FE6
           ,x"ffff" -- 7FE8
           ,x"ffff" -- 7FEA
           ,x"ffff" -- 7FEC
           ,x"ffff" -- 7FEE
           ,x"ffff" -- 7FF0
           ,x"ffff" -- 7FF2
           ,x"ffff" -- 7FF4
           ,x"ffff" -- 7FF6
           ,x"ffff" -- 7FF8
           ,x"ffff" -- 7FFA
           ,x"ffff" -- 7FFC
           ,x"ffff" -- 7FFE
	);
begin

	process(clk)
	variable addr_int : integer range 0 to romLast := 0;
	begin
		if rising_edge(clk) then
			addr_int := to_integer( unsigned( addr ));	-- word address
			data_out <= pgmRom( addr_int );
		end if;
	end process;

end Behavioral;
  